magic
tech gf180mcuD
timestamp 1765407047
<< metal1 >>
rect 2775 2610 2850 2625
rect 2715 2595 2850 2610
rect 2670 2580 2835 2595
rect 2625 2565 2835 2580
rect 2580 2550 2835 2565
rect 2550 2535 2835 2550
rect 1275 2520 1590 2535
rect 2520 2520 2820 2535
rect 1185 2505 1680 2520
rect 2490 2505 2820 2520
rect 1125 2490 1740 2505
rect 2460 2490 2820 2505
rect 1080 2475 1785 2490
rect 2445 2475 2820 2490
rect 1035 2460 1830 2475
rect 2415 2460 2805 2475
rect 1005 2445 1860 2460
rect 2400 2445 2805 2460
rect 975 2430 1890 2445
rect 2370 2430 2805 2445
rect 240 2370 255 2430
rect 945 2415 1395 2430
rect 1470 2415 1920 2430
rect 2355 2415 2790 2430
rect 915 2400 1260 2415
rect 1605 2400 1950 2415
rect 2340 2400 2790 2415
rect 885 2385 1185 2400
rect 1680 2385 1980 2400
rect 2310 2385 2775 2400
rect 855 2370 1125 2385
rect 1740 2370 2010 2385
rect 2295 2370 2775 2385
rect 225 2340 270 2370
rect 840 2355 1080 2370
rect 1785 2355 2040 2370
rect 2280 2355 2775 2370
rect 810 2340 1050 2355
rect 1815 2340 2055 2355
rect 2265 2340 2430 2355
rect 2535 2340 2760 2355
rect 210 2325 285 2340
rect 780 2325 1005 2340
rect 1860 2325 2085 2340
rect 2235 2325 2415 2340
rect 2550 2325 2760 2340
rect 195 2310 285 2325
rect 765 2310 975 2325
rect 1890 2310 2100 2325
rect 2220 2310 2400 2325
rect 180 2295 300 2310
rect 750 2295 945 2310
rect 1920 2295 2115 2310
rect 2205 2295 2400 2310
rect 2565 2295 2745 2325
rect 180 2280 315 2295
rect 720 2280 930 2295
rect 1935 2280 2100 2295
rect 2190 2280 2400 2295
rect 150 2265 330 2280
rect 705 2265 900 2280
rect 1965 2265 2085 2280
rect 2175 2265 2400 2280
rect 2580 2280 2730 2295
rect 2580 2265 2715 2280
rect 135 2250 360 2265
rect 690 2250 870 2265
rect 1995 2250 2070 2265
rect 2160 2250 2400 2265
rect 120 2235 375 2250
rect 675 2235 855 2250
rect 2010 2235 2070 2250
rect 2145 2235 2400 2250
rect 90 2220 405 2235
rect 660 2220 840 2235
rect 2025 2220 2055 2235
rect 2130 2220 2400 2235
rect 2565 2250 2715 2265
rect 2565 2220 2700 2250
rect 15 2205 465 2220
rect 645 2205 810 2220
rect 2115 2205 2415 2220
rect 2550 2205 2685 2220
rect 90 2190 405 2205
rect 630 2190 795 2205
rect 2100 2190 2430 2205
rect 2535 2190 2670 2205
rect 120 2175 375 2190
rect 615 2175 780 2190
rect 2100 2175 2475 2190
rect 2505 2175 2670 2190
rect 135 2160 345 2175
rect 600 2160 765 2175
rect 2085 2160 2655 2175
rect 165 2145 330 2160
rect 585 2145 750 2160
rect 2070 2145 2640 2160
rect 180 2130 315 2145
rect 570 2130 735 2145
rect 2055 2130 2625 2145
rect 195 2115 300 2130
rect 570 2115 720 2130
rect 2040 2115 2625 2130
rect 195 2100 285 2115
rect 555 2100 705 2115
rect 2025 2100 2610 2115
rect 210 2085 285 2100
rect 540 2085 690 2100
rect 1995 2085 2595 2100
rect 225 2055 270 2085
rect 525 2070 675 2085
rect 1845 2070 2580 2085
rect 525 2055 660 2070
rect 1800 2055 2565 2070
rect 240 1995 255 2055
rect 510 2040 645 2055
rect 1785 2040 2565 2055
rect 495 2025 645 2040
rect 1770 2025 2550 2040
rect 495 2010 630 2025
rect 1755 2010 2535 2025
rect 480 1995 615 2010
rect 1725 1995 2520 2010
rect 465 1965 600 1995
rect 1710 1980 2505 1995
rect 1695 1965 2490 1980
rect 450 1950 585 1965
rect 1665 1950 2475 1965
rect 450 1935 570 1950
rect 1650 1935 2460 1950
rect 435 1920 570 1935
rect 1620 1920 2445 1935
rect 435 1905 555 1920
rect 1605 1905 2430 1920
rect 420 1890 555 1905
rect 1590 1890 2415 1905
rect 420 1875 540 1890
rect 1575 1875 2385 1890
rect 405 1860 540 1875
rect 1545 1860 2370 1875
rect 405 1845 525 1860
rect 1530 1845 2355 1860
rect 2445 1845 2460 1860
rect 390 1830 525 1845
rect 1515 1830 2340 1845
rect 2430 1830 2475 1845
rect 390 1800 510 1830
rect 690 1815 735 1830
rect 1020 1815 1080 1830
rect 1350 1815 1410 1830
rect 1665 1815 2325 1830
rect 2415 1815 2475 1830
rect 675 1800 750 1815
rect 1005 1800 1095 1815
rect 1335 1800 1425 1815
rect 375 1755 495 1800
rect 660 1785 765 1800
rect 990 1785 1110 1800
rect 1320 1785 1440 1800
rect 645 1770 780 1785
rect 975 1770 1125 1785
rect 1305 1770 1455 1785
rect 1815 1770 2295 1815
rect 2400 1800 2490 1815
rect 2385 1785 2490 1800
rect 630 1755 705 1770
rect 735 1755 795 1770
rect 960 1755 1035 1770
rect 1065 1755 1140 1770
rect 1290 1755 1365 1770
rect 1395 1755 1470 1770
rect 360 1710 480 1755
rect 615 1740 690 1755
rect 750 1740 810 1755
rect 945 1740 1005 1755
rect 1080 1740 1155 1755
rect 1275 1740 1350 1755
rect 1410 1740 1485 1755
rect 1800 1740 2295 1770
rect 2370 1770 2490 1785
rect 2370 1755 2505 1770
rect 600 1725 675 1740
rect 765 1725 840 1740
rect 930 1725 990 1740
rect 1095 1725 1170 1740
rect 1260 1725 1335 1740
rect 1425 1725 1500 1740
rect 585 1710 660 1725
rect 780 1710 855 1725
rect 915 1710 975 1725
rect 1110 1710 1185 1725
rect 1245 1710 1320 1725
rect 1440 1710 1515 1725
rect 1785 1710 2295 1740
rect 2385 1725 2505 1755
rect 2385 1710 2520 1725
rect 345 1650 465 1710
rect 570 1695 645 1710
rect 795 1695 870 1710
rect 900 1695 960 1710
rect 1125 1695 1200 1710
rect 1230 1695 1305 1710
rect 1455 1695 1530 1710
rect 1800 1695 2295 1710
rect 555 1680 630 1695
rect 810 1680 945 1695
rect 1140 1680 1290 1695
rect 1470 1680 1545 1695
rect 1815 1680 2280 1695
rect 540 1665 600 1680
rect 825 1665 930 1680
rect 1155 1665 1275 1680
rect 1485 1665 1560 1680
rect 1830 1665 2280 1680
rect 2400 1665 2520 1710
rect 525 1650 585 1665
rect 330 1575 450 1650
rect 525 1635 600 1650
rect 840 1635 930 1665
rect 1170 1635 1260 1665
rect 1500 1635 1560 1665
rect 1740 1650 1755 1665
rect 1860 1650 2280 1665
rect 540 1620 600 1635
rect 825 1620 930 1635
rect 1155 1620 1275 1635
rect 1485 1620 1560 1635
rect 1725 1635 1770 1650
rect 1725 1620 1785 1635
rect 1875 1620 2280 1650
rect 555 1605 630 1620
rect 810 1605 945 1620
rect 1140 1605 1290 1620
rect 1470 1605 1545 1620
rect 1710 1605 1800 1620
rect 1890 1605 2010 1620
rect 2025 1605 2280 1620
rect 2415 1650 2520 1665
rect 570 1590 645 1605
rect 795 1590 870 1605
rect 900 1590 960 1605
rect 1125 1590 1200 1605
rect 1230 1590 1305 1605
rect 1455 1590 1530 1605
rect 1695 1590 1815 1605
rect 1905 1590 1965 1605
rect 2025 1590 2265 1605
rect 2415 1590 2535 1650
rect 585 1575 660 1590
rect 780 1575 855 1590
rect 915 1575 975 1590
rect 1110 1575 1185 1590
rect 1245 1575 1320 1590
rect 1440 1575 1515 1590
rect 1680 1575 1830 1590
rect 1920 1575 1935 1590
rect 2025 1575 2250 1590
rect 315 1560 435 1575
rect 600 1560 675 1575
rect 765 1560 840 1575
rect 930 1560 990 1575
rect 1095 1560 1170 1575
rect 1260 1560 1335 1575
rect 1425 1560 1500 1575
rect 1665 1560 1845 1575
rect 300 1530 435 1560
rect 615 1545 690 1560
rect 750 1545 810 1560
rect 945 1545 1005 1560
rect 1080 1545 1155 1560
rect 1275 1545 1350 1560
rect 1410 1545 1485 1560
rect 1650 1545 1860 1560
rect 2025 1545 2235 1575
rect 2430 1560 2535 1590
rect 630 1530 705 1545
rect 735 1530 795 1545
rect 960 1530 1035 1545
rect 1065 1530 1140 1545
rect 1290 1530 1365 1545
rect 1395 1530 1470 1545
rect 1620 1530 1845 1545
rect 2025 1530 2220 1545
rect 285 1515 435 1530
rect 645 1515 780 1530
rect 975 1515 1125 1530
rect 1305 1515 1455 1530
rect 1605 1515 1830 1530
rect 2025 1515 2205 1530
rect 270 1485 435 1515
rect 660 1500 765 1515
rect 990 1500 1110 1515
rect 1320 1500 1440 1515
rect 1590 1500 1815 1515
rect 2025 1500 2190 1515
rect 675 1485 750 1500
rect 255 1455 300 1485
rect 240 1425 285 1455
rect 225 1395 270 1425
rect 210 1380 255 1395
rect 195 1365 255 1380
rect 195 1335 240 1365
rect 180 1320 240 1335
rect 180 1290 225 1320
rect 315 1290 435 1485
rect 690 1470 765 1485
rect 1005 1470 1095 1500
rect 1335 1485 1425 1500
rect 1575 1485 1800 1500
rect 1335 1470 1410 1485
rect 1560 1470 1785 1485
rect 2025 1470 2175 1500
rect 705 1455 780 1470
rect 990 1455 1110 1470
rect 1320 1455 1395 1470
rect 1545 1455 1770 1470
rect 2025 1455 2160 1470
rect 720 1440 795 1455
rect 975 1440 1125 1455
rect 1305 1440 1380 1455
rect 1530 1440 1755 1455
rect 735 1425 795 1440
rect 960 1425 1035 1440
rect 1065 1425 1125 1440
rect 1290 1425 1365 1440
rect 1515 1425 1740 1440
rect 2025 1425 2145 1455
rect 750 1410 810 1425
rect 945 1410 1020 1425
rect 1080 1410 1140 1425
rect 1275 1410 1350 1425
rect 1500 1410 1725 1425
rect 2025 1410 2130 1425
rect 765 1395 840 1410
rect 930 1395 1005 1410
rect 1095 1395 1155 1410
rect 1260 1395 1335 1410
rect 1470 1395 1695 1410
rect 1785 1395 1815 1410
rect 2025 1395 2115 1410
rect 780 1380 855 1395
rect 915 1380 990 1395
rect 1110 1380 1170 1395
rect 1245 1380 1320 1395
rect 1455 1380 1680 1395
rect 1770 1380 1830 1395
rect 795 1365 870 1380
rect 900 1365 975 1380
rect 1125 1365 1185 1380
rect 1230 1365 1305 1380
rect 1440 1365 1665 1380
rect 1755 1365 1845 1380
rect 2025 1365 2100 1395
rect 810 1350 960 1365
rect 1140 1350 1290 1365
rect 1410 1350 1650 1365
rect 1740 1350 1860 1365
rect 2025 1350 2085 1365
rect 825 1335 945 1350
rect 1155 1335 1275 1350
rect 1395 1335 1620 1350
rect 1725 1335 1785 1350
rect 1800 1335 1875 1350
rect 2025 1335 2070 1350
rect 840 1320 930 1335
rect 1170 1320 1260 1335
rect 1380 1320 1605 1335
rect 1710 1320 1770 1335
rect 1815 1320 1890 1335
rect 2025 1320 2055 1335
rect 855 1305 915 1320
rect 1185 1305 1245 1320
rect 1350 1305 1590 1320
rect 1695 1305 1755 1320
rect 1830 1305 1905 1320
rect 2025 1305 2040 1320
rect 870 1290 885 1305
rect 1200 1290 1215 1305
rect 1335 1290 1560 1305
rect 1680 1290 1740 1305
rect 1860 1290 1920 1305
rect 165 1230 225 1290
rect 330 1260 435 1290
rect 1305 1275 1545 1290
rect 1665 1275 1725 1290
rect 1875 1275 1935 1290
rect 2430 1275 2550 1560
rect 1290 1260 1515 1275
rect 1650 1260 1710 1275
rect 1890 1260 1950 1275
rect 165 1170 210 1230
rect 330 1200 450 1260
rect 1260 1245 1500 1260
rect 1620 1245 1695 1260
rect 1905 1245 1965 1260
rect 2430 1245 2535 1275
rect 1245 1230 1470 1245
rect 1605 1230 1680 1245
rect 1215 1215 1455 1230
rect 1605 1215 1665 1230
rect 1200 1200 1440 1215
rect 1590 1200 1680 1215
rect 1920 1200 1980 1245
rect 345 1185 450 1200
rect 1170 1185 1410 1200
rect 1575 1185 1695 1200
rect 1905 1185 1965 1200
rect 2415 1185 2535 1245
rect 165 1110 225 1170
rect 345 1140 465 1185
rect 1155 1170 1380 1185
rect 1560 1170 1620 1185
rect 1635 1170 1710 1185
rect 1890 1170 1950 1185
rect 2415 1170 2520 1185
rect 1125 1155 1365 1170
rect 1545 1155 1605 1170
rect 1650 1155 1725 1170
rect 1875 1155 1935 1170
rect 1095 1140 1335 1155
rect 1530 1140 1590 1155
rect 1665 1140 1740 1155
rect 1860 1140 1920 1155
rect 360 1125 465 1140
rect 1080 1125 1305 1140
rect 1515 1125 1575 1140
rect 1680 1125 1755 1140
rect 1830 1125 1905 1140
rect 2400 1125 2520 1170
rect 165 1095 240 1110
rect 180 1080 240 1095
rect 360 1080 480 1125
rect 1050 1110 1275 1125
rect 1500 1110 1560 1125
rect 1695 1110 1770 1125
rect 1815 1110 1890 1125
rect 1020 1095 1260 1110
rect 1485 1095 1545 1110
rect 1710 1095 1785 1110
rect 1800 1095 1875 1110
rect 990 1080 1230 1095
rect 1470 1080 1530 1095
rect 1725 1080 1860 1095
rect 2385 1080 2505 1125
rect 180 1065 255 1080
rect 180 1050 270 1065
rect 195 1035 270 1050
rect 375 1050 495 1080
rect 960 1065 1200 1080
rect 1455 1065 1515 1080
rect 1740 1065 1845 1080
rect 930 1050 1170 1065
rect 1440 1050 1500 1065
rect 1755 1050 1830 1065
rect 375 1035 510 1050
rect 900 1035 1140 1050
rect 1440 1035 1515 1050
rect 1740 1035 1845 1050
rect 2370 1035 2490 1080
rect 210 1020 300 1035
rect 420 1020 510 1035
rect 855 1020 1110 1035
rect 1455 1020 1530 1035
rect 1725 1020 1860 1035
rect 210 1005 315 1020
rect 480 1005 510 1020
rect 825 1005 1080 1020
rect 1470 1005 1545 1020
rect 1725 1005 1785 1020
rect 1800 1005 1875 1020
rect 2355 1005 2475 1035
rect 225 990 330 1005
rect 780 990 1050 1005
rect 1485 990 1560 1005
rect 1710 990 1770 1005
rect 1815 990 1890 1005
rect 2340 990 2475 1005
rect 240 975 360 990
rect 735 975 1020 990
rect 1500 975 1575 990
rect 1695 975 1755 990
rect 1830 975 1905 990
rect 2340 975 2460 990
rect 255 960 405 975
rect 690 960 975 975
rect 1515 960 1590 975
rect 1680 960 1740 975
rect 1845 960 1920 975
rect 2325 960 2460 975
rect 285 945 480 960
rect 600 945 945 960
rect 1530 945 1605 960
rect 1665 945 1725 960
rect 1860 945 1935 960
rect 2325 945 2445 960
rect 300 930 900 945
rect 1545 930 1620 945
rect 1650 930 1710 945
rect 1875 930 1950 945
rect 2310 930 2445 945
rect 330 915 855 930
rect 1560 915 1695 930
rect 1890 915 1965 930
rect 2310 915 2430 930
rect 360 900 810 915
rect 1575 900 1680 915
rect 1905 900 1980 915
rect 390 885 750 900
rect 1590 885 1665 900
rect 465 870 675 885
rect 1590 870 1680 885
rect 1920 870 1980 900
rect 2295 900 2430 915
rect 2295 885 2415 900
rect 2280 870 2415 885
rect 1575 855 1695 870
rect 1905 855 1965 870
rect 1560 840 1620 855
rect 1635 840 1710 855
rect 1890 840 1950 855
rect 2265 840 2400 870
rect 2640 855 2655 870
rect 2625 840 2655 855
rect 1545 825 1605 840
rect 1650 825 1725 840
rect 1875 825 1935 840
rect 2250 825 2385 840
rect 1530 810 1590 825
rect 1665 810 1740 825
rect 1860 810 1920 825
rect 2235 810 2370 825
rect 2625 810 2670 840
rect 495 795 645 810
rect 1515 795 1575 810
rect 1680 795 1755 810
rect 1845 795 1905 810
rect 2220 795 2370 810
rect 2610 795 2685 810
rect 510 780 660 795
rect 1500 780 1560 795
rect 1695 780 1770 795
rect 1830 780 1890 795
rect 2220 780 2355 795
rect 2595 780 2700 795
rect 525 765 660 780
rect 1485 765 1545 780
rect 1710 765 1785 780
rect 1815 765 1875 780
rect 2205 765 2340 780
rect 2580 765 2715 780
rect 525 750 675 765
rect 1470 750 1530 765
rect 1725 750 1860 765
rect 2190 750 2340 765
rect 2550 750 2745 765
rect 540 735 690 750
rect 1455 735 1515 750
rect 1740 735 1845 750
rect 2175 735 2325 750
rect 2520 735 2775 750
rect 555 720 705 735
rect 1440 720 1500 735
rect 1755 720 1830 735
rect 2160 720 2310 735
rect 2565 720 2730 735
rect 570 705 720 720
rect 1440 705 1515 720
rect 1755 705 1815 720
rect 2145 705 2295 720
rect 2580 705 2700 720
rect 585 690 735 705
rect 1455 690 1530 705
rect 1740 690 1800 705
rect 2130 690 2295 705
rect 2595 690 2685 705
rect 600 675 750 690
rect 1470 675 1545 690
rect 1725 675 1785 690
rect 2115 675 2280 690
rect 2610 675 2670 690
rect 600 660 765 675
rect 1485 660 1560 675
rect 1710 660 1770 675
rect 2100 660 2265 675
rect 2625 660 2670 675
rect 630 645 780 660
rect 1500 645 1575 660
rect 1695 645 1755 660
rect 2085 645 2250 660
rect 2625 645 2655 660
rect 645 630 810 645
rect 1515 630 1590 645
rect 1680 630 1740 645
rect 2070 630 2235 645
rect 2640 630 2655 645
rect 660 615 825 630
rect 1530 615 1605 630
rect 1665 615 1725 630
rect 2040 615 2220 630
rect 660 600 840 615
rect 1545 600 1605 615
rect 1650 600 1710 615
rect 2025 600 2205 615
rect 675 585 870 600
rect 1560 585 1695 600
rect 2010 585 2190 600
rect 705 570 885 585
rect 1575 570 1680 585
rect 1980 570 2175 585
rect 720 555 915 570
rect 1590 555 1665 570
rect 1965 555 2145 570
rect 735 540 930 555
rect 1605 540 1650 555
rect 1935 540 2130 555
rect 750 525 960 540
rect 1905 525 2115 540
rect 780 510 990 525
rect 1875 510 2100 525
rect 795 495 1020 510
rect 1845 495 2070 510
rect 810 480 1065 495
rect 1800 480 2055 495
rect 840 465 1095 480
rect 1770 465 2025 480
rect 870 450 1155 465
rect 1725 450 1995 465
rect 900 435 1200 450
rect 1665 435 1980 450
rect 915 420 1290 435
rect 1575 420 1950 435
rect 945 405 1920 420
rect 975 390 1890 405
rect 1005 375 1860 390
rect 1050 360 1815 375
rect 1095 345 1770 360
rect 1155 330 1710 345
rect 1215 315 1650 330
rect 1320 300 1545 315
<< metal2 >>
rect 2775 2610 2850 2625
rect 2715 2595 2850 2610
rect 2670 2580 2835 2595
rect 2625 2565 2835 2580
rect 2580 2550 2835 2565
rect 2550 2535 2835 2550
rect 1275 2520 1590 2535
rect 2520 2520 2820 2535
rect 1185 2505 1680 2520
rect 2490 2505 2820 2520
rect 1125 2490 1740 2505
rect 2460 2490 2820 2505
rect 1080 2475 1785 2490
rect 2445 2475 2820 2490
rect 1035 2460 1830 2475
rect 2415 2460 2805 2475
rect 1005 2445 1860 2460
rect 2400 2445 2805 2460
rect 975 2430 1890 2445
rect 2370 2430 2805 2445
rect 240 2370 255 2430
rect 945 2415 1395 2430
rect 1470 2415 1920 2430
rect 2355 2415 2790 2430
rect 915 2400 1260 2415
rect 1605 2400 1950 2415
rect 2340 2400 2790 2415
rect 885 2385 1185 2400
rect 1680 2385 1980 2400
rect 2310 2385 2775 2400
rect 855 2370 1125 2385
rect 1740 2370 2010 2385
rect 2295 2370 2775 2385
rect 225 2340 270 2370
rect 840 2355 1080 2370
rect 1785 2355 2040 2370
rect 2280 2355 2775 2370
rect 810 2340 1050 2355
rect 1815 2340 2055 2355
rect 2265 2340 2430 2355
rect 2535 2340 2760 2355
rect 210 2325 285 2340
rect 780 2325 1005 2340
rect 1860 2325 2085 2340
rect 2235 2325 2415 2340
rect 2550 2325 2760 2340
rect 195 2310 285 2325
rect 765 2310 975 2325
rect 1890 2310 2100 2325
rect 2220 2310 2400 2325
rect 180 2295 300 2310
rect 750 2295 945 2310
rect 1920 2295 2115 2310
rect 2205 2295 2400 2310
rect 2565 2295 2745 2325
rect 180 2280 315 2295
rect 720 2280 930 2295
rect 1935 2280 2100 2295
rect 2190 2280 2400 2295
rect 150 2265 330 2280
rect 705 2265 900 2280
rect 1965 2265 2085 2280
rect 2175 2265 2400 2280
rect 2580 2280 2730 2295
rect 2580 2265 2715 2280
rect 135 2250 360 2265
rect 690 2250 870 2265
rect 1995 2250 2070 2265
rect 2160 2250 2400 2265
rect 120 2235 375 2250
rect 675 2235 855 2250
rect 2010 2235 2070 2250
rect 2145 2235 2400 2250
rect 90 2220 405 2235
rect 660 2220 840 2235
rect 2025 2220 2055 2235
rect 2130 2220 2400 2235
rect 2565 2250 2715 2265
rect 2565 2220 2700 2250
rect 15 2205 465 2220
rect 645 2205 810 2220
rect 2115 2205 2415 2220
rect 2550 2205 2685 2220
rect 90 2190 405 2205
rect 630 2190 795 2205
rect 2100 2190 2430 2205
rect 2535 2190 2670 2205
rect 120 2175 375 2190
rect 615 2175 780 2190
rect 2100 2175 2475 2190
rect 2505 2175 2670 2190
rect 135 2160 345 2175
rect 600 2160 765 2175
rect 2085 2160 2655 2175
rect 165 2145 330 2160
rect 585 2145 750 2160
rect 2070 2145 2640 2160
rect 180 2130 315 2145
rect 570 2130 735 2145
rect 2055 2130 2625 2145
rect 195 2115 300 2130
rect 570 2115 720 2130
rect 2040 2115 2625 2130
rect 195 2100 285 2115
rect 555 2100 705 2115
rect 2025 2100 2610 2115
rect 210 2085 285 2100
rect 540 2085 690 2100
rect 1995 2085 2595 2100
rect 225 2055 270 2085
rect 525 2070 675 2085
rect 1845 2070 2580 2085
rect 525 2055 660 2070
rect 1800 2055 2565 2070
rect 240 1995 255 2055
rect 510 2040 645 2055
rect 1785 2040 2565 2055
rect 495 2025 645 2040
rect 1770 2025 2550 2040
rect 495 2010 630 2025
rect 1755 2010 2535 2025
rect 480 1995 615 2010
rect 1725 1995 2520 2010
rect 465 1965 600 1995
rect 1710 1980 2505 1995
rect 1695 1965 2490 1980
rect 450 1950 585 1965
rect 1665 1950 2475 1965
rect 450 1935 570 1950
rect 1650 1935 2460 1950
rect 435 1920 570 1935
rect 1620 1920 2445 1935
rect 435 1905 555 1920
rect 1605 1905 2430 1920
rect 420 1890 555 1905
rect 1590 1890 2415 1905
rect 420 1875 540 1890
rect 1575 1875 2385 1890
rect 405 1860 540 1875
rect 1545 1860 2370 1875
rect 405 1845 525 1860
rect 1530 1845 2355 1860
rect 2445 1845 2460 1860
rect 390 1830 525 1845
rect 1515 1830 2340 1845
rect 2430 1830 2475 1845
rect 390 1800 510 1830
rect 690 1815 735 1830
rect 1020 1815 1080 1830
rect 1350 1815 1410 1830
rect 1665 1815 2325 1830
rect 2415 1815 2475 1830
rect 675 1800 750 1815
rect 1005 1800 1095 1815
rect 1335 1800 1425 1815
rect 375 1755 495 1800
rect 660 1785 765 1800
rect 990 1785 1110 1800
rect 1320 1785 1440 1800
rect 645 1770 780 1785
rect 975 1770 1125 1785
rect 1305 1770 1455 1785
rect 1815 1770 2295 1815
rect 2400 1800 2490 1815
rect 2385 1785 2490 1800
rect 630 1755 705 1770
rect 735 1755 795 1770
rect 960 1755 1035 1770
rect 1065 1755 1140 1770
rect 1290 1755 1365 1770
rect 1395 1755 1470 1770
rect 360 1710 480 1755
rect 615 1740 690 1755
rect 750 1740 810 1755
rect 945 1740 1005 1755
rect 1080 1740 1155 1755
rect 1275 1740 1350 1755
rect 1410 1740 1485 1755
rect 1800 1740 2295 1770
rect 2370 1770 2490 1785
rect 2370 1755 2505 1770
rect 600 1725 675 1740
rect 765 1725 840 1740
rect 930 1725 990 1740
rect 1095 1725 1170 1740
rect 1260 1725 1335 1740
rect 1425 1725 1500 1740
rect 585 1710 660 1725
rect 780 1710 855 1725
rect 915 1710 975 1725
rect 1110 1710 1185 1725
rect 1245 1710 1320 1725
rect 1440 1710 1515 1725
rect 1785 1710 2295 1740
rect 2385 1725 2505 1755
rect 2385 1710 2520 1725
rect 345 1650 465 1710
rect 570 1695 645 1710
rect 795 1695 870 1710
rect 900 1695 960 1710
rect 1125 1695 1200 1710
rect 1230 1695 1305 1710
rect 1455 1695 1530 1710
rect 1800 1695 2295 1710
rect 555 1680 630 1695
rect 810 1680 945 1695
rect 1140 1680 1290 1695
rect 1470 1680 1545 1695
rect 1815 1680 2280 1695
rect 540 1665 600 1680
rect 825 1665 930 1680
rect 1155 1665 1275 1680
rect 1485 1665 1560 1680
rect 1830 1665 2280 1680
rect 2400 1665 2520 1710
rect 525 1650 585 1665
rect 330 1575 450 1650
rect 525 1635 600 1650
rect 840 1635 930 1665
rect 1170 1635 1260 1665
rect 1500 1635 1560 1665
rect 1740 1650 1755 1665
rect 1860 1650 2280 1665
rect 540 1620 600 1635
rect 825 1620 930 1635
rect 1155 1620 1275 1635
rect 1485 1620 1560 1635
rect 1725 1635 1770 1650
rect 1725 1620 1785 1635
rect 1875 1620 2280 1650
rect 555 1605 630 1620
rect 810 1605 945 1620
rect 1140 1605 1290 1620
rect 1470 1605 1545 1620
rect 1710 1605 1800 1620
rect 1890 1605 2010 1620
rect 2025 1605 2280 1620
rect 2415 1650 2520 1665
rect 570 1590 645 1605
rect 795 1590 870 1605
rect 900 1590 960 1605
rect 1125 1590 1200 1605
rect 1230 1590 1305 1605
rect 1455 1590 1530 1605
rect 1695 1590 1815 1605
rect 1905 1590 1965 1605
rect 2025 1590 2265 1605
rect 2415 1590 2535 1650
rect 585 1575 660 1590
rect 780 1575 855 1590
rect 915 1575 975 1590
rect 1110 1575 1185 1590
rect 1245 1575 1320 1590
rect 1440 1575 1515 1590
rect 1680 1575 1830 1590
rect 1920 1575 1935 1590
rect 2025 1575 2250 1590
rect 315 1560 435 1575
rect 600 1560 675 1575
rect 765 1560 840 1575
rect 930 1560 990 1575
rect 1095 1560 1170 1575
rect 1260 1560 1335 1575
rect 1425 1560 1500 1575
rect 1665 1560 1845 1575
rect 300 1530 435 1560
rect 615 1545 690 1560
rect 750 1545 810 1560
rect 945 1545 1005 1560
rect 1080 1545 1155 1560
rect 1275 1545 1350 1560
rect 1410 1545 1485 1560
rect 1650 1545 1860 1560
rect 2025 1545 2235 1575
rect 2430 1560 2535 1590
rect 630 1530 705 1545
rect 735 1530 795 1545
rect 960 1530 1035 1545
rect 1065 1530 1140 1545
rect 1290 1530 1365 1545
rect 1395 1530 1470 1545
rect 1620 1530 1845 1545
rect 2025 1530 2220 1545
rect 285 1515 435 1530
rect 645 1515 780 1530
rect 975 1515 1125 1530
rect 1305 1515 1455 1530
rect 1605 1515 1830 1530
rect 2025 1515 2205 1530
rect 270 1485 435 1515
rect 660 1500 765 1515
rect 990 1500 1110 1515
rect 1320 1500 1440 1515
rect 1590 1500 1815 1515
rect 2025 1500 2190 1515
rect 675 1485 750 1500
rect 255 1455 300 1485
rect 240 1425 285 1455
rect 225 1395 270 1425
rect 210 1380 255 1395
rect 195 1365 255 1380
rect 195 1335 240 1365
rect 180 1320 240 1335
rect 180 1290 225 1320
rect 315 1290 435 1485
rect 690 1470 765 1485
rect 1005 1470 1095 1500
rect 1335 1485 1425 1500
rect 1575 1485 1800 1500
rect 1335 1470 1410 1485
rect 1560 1470 1785 1485
rect 2025 1470 2175 1500
rect 705 1455 780 1470
rect 990 1455 1110 1470
rect 1320 1455 1395 1470
rect 1545 1455 1770 1470
rect 2025 1455 2160 1470
rect 720 1440 795 1455
rect 975 1440 1125 1455
rect 1305 1440 1380 1455
rect 1530 1440 1755 1455
rect 735 1425 795 1440
rect 960 1425 1035 1440
rect 1065 1425 1125 1440
rect 1290 1425 1365 1440
rect 1515 1425 1740 1440
rect 2025 1425 2145 1455
rect 750 1410 810 1425
rect 945 1410 1020 1425
rect 1080 1410 1140 1425
rect 1275 1410 1350 1425
rect 1500 1410 1725 1425
rect 2025 1410 2130 1425
rect 765 1395 840 1410
rect 930 1395 1005 1410
rect 1095 1395 1155 1410
rect 1260 1395 1335 1410
rect 1470 1395 1695 1410
rect 1785 1395 1815 1410
rect 2025 1395 2115 1410
rect 780 1380 855 1395
rect 915 1380 990 1395
rect 1110 1380 1170 1395
rect 1245 1380 1320 1395
rect 1455 1380 1680 1395
rect 1770 1380 1830 1395
rect 795 1365 870 1380
rect 900 1365 975 1380
rect 1125 1365 1185 1380
rect 1230 1365 1305 1380
rect 1440 1365 1665 1380
rect 1755 1365 1845 1380
rect 2025 1365 2100 1395
rect 810 1350 960 1365
rect 1140 1350 1290 1365
rect 1410 1350 1650 1365
rect 1740 1350 1860 1365
rect 2025 1350 2085 1365
rect 825 1335 945 1350
rect 1155 1335 1275 1350
rect 1395 1335 1620 1350
rect 1725 1335 1785 1350
rect 1800 1335 1875 1350
rect 2025 1335 2070 1350
rect 840 1320 930 1335
rect 1170 1320 1260 1335
rect 1380 1320 1605 1335
rect 1710 1320 1770 1335
rect 1815 1320 1890 1335
rect 2025 1320 2055 1335
rect 855 1305 915 1320
rect 1185 1305 1245 1320
rect 1350 1305 1590 1320
rect 1695 1305 1755 1320
rect 1830 1305 1905 1320
rect 2025 1305 2040 1320
rect 870 1290 885 1305
rect 1200 1290 1215 1305
rect 1335 1290 1560 1305
rect 1680 1290 1740 1305
rect 1860 1290 1920 1305
rect 165 1230 225 1290
rect 330 1260 435 1290
rect 1305 1275 1545 1290
rect 1665 1275 1725 1290
rect 1875 1275 1935 1290
rect 2430 1275 2550 1560
rect 1290 1260 1515 1275
rect 1650 1260 1710 1275
rect 1890 1260 1950 1275
rect 165 1170 210 1230
rect 330 1200 450 1260
rect 1260 1245 1500 1260
rect 1620 1245 1695 1260
rect 1905 1245 1965 1260
rect 2430 1245 2535 1275
rect 1245 1230 1470 1245
rect 1605 1230 1680 1245
rect 1215 1215 1455 1230
rect 1605 1215 1665 1230
rect 1200 1200 1440 1215
rect 1590 1200 1680 1215
rect 1920 1200 1980 1245
rect 345 1185 450 1200
rect 1170 1185 1410 1200
rect 1575 1185 1695 1200
rect 1905 1185 1965 1200
rect 2415 1185 2535 1245
rect 165 1110 225 1170
rect 345 1140 465 1185
rect 1155 1170 1380 1185
rect 1560 1170 1620 1185
rect 1635 1170 1710 1185
rect 1890 1170 1950 1185
rect 2415 1170 2520 1185
rect 1125 1155 1365 1170
rect 1545 1155 1605 1170
rect 1650 1155 1725 1170
rect 1875 1155 1935 1170
rect 1095 1140 1335 1155
rect 1530 1140 1590 1155
rect 1665 1140 1740 1155
rect 1860 1140 1920 1155
rect 360 1125 465 1140
rect 1080 1125 1305 1140
rect 1515 1125 1575 1140
rect 1680 1125 1755 1140
rect 1830 1125 1905 1140
rect 2400 1125 2520 1170
rect 165 1095 240 1110
rect 180 1080 240 1095
rect 360 1080 480 1125
rect 1050 1110 1275 1125
rect 1500 1110 1560 1125
rect 1695 1110 1770 1125
rect 1815 1110 1890 1125
rect 1020 1095 1260 1110
rect 1485 1095 1545 1110
rect 1710 1095 1785 1110
rect 1800 1095 1875 1110
rect 990 1080 1230 1095
rect 1470 1080 1530 1095
rect 1725 1080 1860 1095
rect 2385 1080 2505 1125
rect 180 1065 255 1080
rect 180 1050 270 1065
rect 195 1035 270 1050
rect 375 1050 495 1080
rect 960 1065 1200 1080
rect 1455 1065 1515 1080
rect 1740 1065 1845 1080
rect 930 1050 1170 1065
rect 1440 1050 1500 1065
rect 1755 1050 1830 1065
rect 375 1035 510 1050
rect 900 1035 1140 1050
rect 1440 1035 1515 1050
rect 1740 1035 1845 1050
rect 2370 1035 2490 1080
rect 210 1020 300 1035
rect 420 1020 510 1035
rect 855 1020 1110 1035
rect 1455 1020 1530 1035
rect 1725 1020 1860 1035
rect 210 1005 315 1020
rect 480 1005 510 1020
rect 825 1005 1080 1020
rect 1470 1005 1545 1020
rect 1725 1005 1785 1020
rect 1800 1005 1875 1020
rect 2355 1005 2475 1035
rect 225 990 330 1005
rect 780 990 1050 1005
rect 1485 990 1560 1005
rect 1710 990 1770 1005
rect 1815 990 1890 1005
rect 2340 990 2475 1005
rect 240 975 360 990
rect 735 975 1020 990
rect 1500 975 1575 990
rect 1695 975 1755 990
rect 1830 975 1905 990
rect 2340 975 2460 990
rect 255 960 405 975
rect 690 960 975 975
rect 1515 960 1590 975
rect 1680 960 1740 975
rect 1845 960 1920 975
rect 2325 960 2460 975
rect 285 945 480 960
rect 600 945 945 960
rect 1530 945 1605 960
rect 1665 945 1725 960
rect 1860 945 1935 960
rect 2325 945 2445 960
rect 300 930 900 945
rect 1545 930 1620 945
rect 1650 930 1710 945
rect 1875 930 1950 945
rect 2310 930 2445 945
rect 330 915 855 930
rect 1560 915 1695 930
rect 1890 915 1965 930
rect 2310 915 2430 930
rect 360 900 810 915
rect 1575 900 1680 915
rect 1905 900 1980 915
rect 390 885 750 900
rect 1590 885 1665 900
rect 465 870 675 885
rect 1590 870 1680 885
rect 1920 870 1980 900
rect 2295 900 2430 915
rect 2295 885 2415 900
rect 2280 870 2415 885
rect 1575 855 1695 870
rect 1905 855 1965 870
rect 1560 840 1620 855
rect 1635 840 1710 855
rect 1890 840 1950 855
rect 2265 840 2400 870
rect 2640 855 2655 870
rect 2625 840 2655 855
rect 1545 825 1605 840
rect 1650 825 1725 840
rect 1875 825 1935 840
rect 2250 825 2385 840
rect 1530 810 1590 825
rect 1665 810 1740 825
rect 1860 810 1920 825
rect 2235 810 2370 825
rect 2625 810 2670 840
rect 495 795 645 810
rect 1515 795 1575 810
rect 1680 795 1755 810
rect 1845 795 1905 810
rect 2220 795 2370 810
rect 2610 795 2685 810
rect 510 780 660 795
rect 1500 780 1560 795
rect 1695 780 1770 795
rect 1830 780 1890 795
rect 2220 780 2355 795
rect 2595 780 2700 795
rect 525 765 660 780
rect 1485 765 1545 780
rect 1710 765 1785 780
rect 1815 765 1875 780
rect 2205 765 2340 780
rect 2580 765 2715 780
rect 525 750 675 765
rect 1470 750 1530 765
rect 1725 750 1860 765
rect 2190 750 2340 765
rect 2550 750 2745 765
rect 540 735 690 750
rect 1455 735 1515 750
rect 1740 735 1845 750
rect 2175 735 2325 750
rect 2520 735 2775 750
rect 555 720 705 735
rect 1440 720 1500 735
rect 1755 720 1830 735
rect 2160 720 2310 735
rect 2565 720 2730 735
rect 570 705 720 720
rect 1440 705 1515 720
rect 1755 705 1815 720
rect 2145 705 2295 720
rect 2580 705 2700 720
rect 585 690 735 705
rect 1455 690 1530 705
rect 1740 690 1800 705
rect 2130 690 2295 705
rect 2595 690 2685 705
rect 600 675 750 690
rect 1470 675 1545 690
rect 1725 675 1785 690
rect 2115 675 2280 690
rect 2610 675 2670 690
rect 600 660 765 675
rect 1485 660 1560 675
rect 1710 660 1770 675
rect 2100 660 2265 675
rect 2625 660 2670 675
rect 630 645 780 660
rect 1500 645 1575 660
rect 1695 645 1755 660
rect 2085 645 2250 660
rect 2625 645 2655 660
rect 645 630 810 645
rect 1515 630 1590 645
rect 1680 630 1740 645
rect 2070 630 2235 645
rect 2640 630 2655 645
rect 660 615 825 630
rect 1530 615 1605 630
rect 1665 615 1725 630
rect 2040 615 2220 630
rect 660 600 840 615
rect 1545 600 1605 615
rect 1650 600 1710 615
rect 2025 600 2205 615
rect 675 585 870 600
rect 1560 585 1695 600
rect 2010 585 2190 600
rect 705 570 885 585
rect 1575 570 1680 585
rect 1980 570 2175 585
rect 720 555 915 570
rect 1590 555 1665 570
rect 1965 555 2145 570
rect 735 540 930 555
rect 1605 540 1650 555
rect 1935 540 2130 555
rect 750 525 960 540
rect 1905 525 2115 540
rect 780 510 990 525
rect 1875 510 2100 525
rect 795 495 1020 510
rect 1845 495 2070 510
rect 810 480 1065 495
rect 1800 480 2055 495
rect 840 465 1095 480
rect 1770 465 2025 480
rect 870 450 1155 465
rect 1725 450 1995 465
rect 900 435 1200 450
rect 1665 435 1980 450
rect 915 420 1290 435
rect 1575 420 1950 435
rect 945 405 1920 420
rect 975 390 1890 405
rect 1005 375 1860 390
rect 1050 360 1815 375
rect 1095 345 1770 360
rect 1155 330 1710 345
rect 1215 315 1650 330
rect 1320 300 1545 315
<< metal3 >>
rect 2775 2610 2850 2625
rect 2715 2595 2850 2610
rect 2670 2580 2835 2595
rect 2625 2565 2835 2580
rect 2580 2550 2835 2565
rect 2550 2535 2835 2550
rect 1275 2520 1590 2535
rect 2520 2520 2820 2535
rect 1185 2505 1680 2520
rect 2490 2505 2820 2520
rect 1125 2490 1740 2505
rect 2460 2490 2820 2505
rect 1080 2475 1785 2490
rect 2445 2475 2820 2490
rect 1035 2460 1830 2475
rect 2415 2460 2805 2475
rect 1005 2445 1860 2460
rect 2400 2445 2805 2460
rect 975 2430 1890 2445
rect 2370 2430 2805 2445
rect 240 2370 255 2430
rect 945 2415 1395 2430
rect 1470 2415 1920 2430
rect 2355 2415 2790 2430
rect 915 2400 1260 2415
rect 1605 2400 1950 2415
rect 2340 2400 2790 2415
rect 885 2385 1185 2400
rect 1680 2385 1980 2400
rect 2310 2385 2775 2400
rect 855 2370 1125 2385
rect 1740 2370 2010 2385
rect 2295 2370 2775 2385
rect 225 2340 270 2370
rect 840 2355 1080 2370
rect 1785 2355 2040 2370
rect 2280 2355 2775 2370
rect 810 2340 1050 2355
rect 1815 2340 2055 2355
rect 2265 2340 2430 2355
rect 2535 2340 2760 2355
rect 210 2325 285 2340
rect 780 2325 1005 2340
rect 1860 2325 2085 2340
rect 2235 2325 2415 2340
rect 2550 2325 2760 2340
rect 195 2310 285 2325
rect 765 2310 975 2325
rect 1890 2310 2100 2325
rect 2220 2310 2400 2325
rect 180 2295 300 2310
rect 750 2295 945 2310
rect 1920 2295 2115 2310
rect 2205 2295 2400 2310
rect 2565 2295 2745 2325
rect 180 2280 315 2295
rect 720 2280 930 2295
rect 1935 2280 2100 2295
rect 2190 2280 2400 2295
rect 150 2265 330 2280
rect 705 2265 900 2280
rect 1965 2265 2085 2280
rect 2175 2265 2400 2280
rect 2580 2280 2730 2295
rect 2580 2265 2715 2280
rect 135 2250 360 2265
rect 690 2250 870 2265
rect 1995 2250 2070 2265
rect 2160 2250 2400 2265
rect 120 2235 375 2250
rect 675 2235 855 2250
rect 2010 2235 2070 2250
rect 2145 2235 2400 2250
rect 90 2220 405 2235
rect 660 2220 840 2235
rect 2025 2220 2055 2235
rect 2130 2220 2400 2235
rect 2565 2250 2715 2265
rect 2565 2220 2700 2250
rect 15 2205 465 2220
rect 645 2205 810 2220
rect 2115 2205 2415 2220
rect 2550 2205 2685 2220
rect 90 2190 405 2205
rect 630 2190 795 2205
rect 2100 2190 2430 2205
rect 2535 2190 2670 2205
rect 120 2175 375 2190
rect 615 2175 780 2190
rect 2100 2175 2475 2190
rect 2505 2175 2670 2190
rect 135 2160 345 2175
rect 600 2160 765 2175
rect 2085 2160 2655 2175
rect 165 2145 330 2160
rect 585 2145 750 2160
rect 2070 2145 2640 2160
rect 180 2130 315 2145
rect 570 2130 735 2145
rect 2055 2130 2625 2145
rect 195 2115 300 2130
rect 570 2115 720 2130
rect 2040 2115 2625 2130
rect 195 2100 285 2115
rect 555 2100 705 2115
rect 2025 2100 2610 2115
rect 210 2085 285 2100
rect 540 2085 690 2100
rect 1995 2085 2595 2100
rect 225 2055 270 2085
rect 525 2070 675 2085
rect 1845 2070 2580 2085
rect 525 2055 660 2070
rect 1800 2055 2565 2070
rect 240 1995 255 2055
rect 510 2040 645 2055
rect 1785 2040 2565 2055
rect 495 2025 645 2040
rect 1770 2025 2550 2040
rect 495 2010 630 2025
rect 1755 2010 2535 2025
rect 480 1995 615 2010
rect 1725 1995 2520 2010
rect 465 1965 600 1995
rect 1710 1980 2505 1995
rect 1695 1965 2490 1980
rect 450 1950 585 1965
rect 1665 1950 2475 1965
rect 450 1935 570 1950
rect 1650 1935 2460 1950
rect 435 1920 570 1935
rect 1620 1920 2445 1935
rect 435 1905 555 1920
rect 1605 1905 2430 1920
rect 420 1890 555 1905
rect 1590 1890 2415 1905
rect 420 1875 540 1890
rect 1575 1875 2385 1890
rect 405 1860 540 1875
rect 1545 1860 2370 1875
rect 405 1845 525 1860
rect 1530 1845 2355 1860
rect 2445 1845 2460 1860
rect 390 1830 525 1845
rect 1515 1830 2340 1845
rect 2430 1830 2475 1845
rect 390 1800 510 1830
rect 690 1815 735 1830
rect 1020 1815 1080 1830
rect 1350 1815 1410 1830
rect 1665 1815 2325 1830
rect 2415 1815 2475 1830
rect 675 1800 750 1815
rect 1005 1800 1095 1815
rect 1335 1800 1425 1815
rect 375 1755 495 1800
rect 660 1785 765 1800
rect 990 1785 1110 1800
rect 1320 1785 1440 1800
rect 645 1770 780 1785
rect 975 1770 1125 1785
rect 1305 1770 1455 1785
rect 1815 1770 2295 1815
rect 2400 1800 2490 1815
rect 2385 1785 2490 1800
rect 630 1755 705 1770
rect 735 1755 795 1770
rect 960 1755 1035 1770
rect 1065 1755 1140 1770
rect 1290 1755 1365 1770
rect 1395 1755 1470 1770
rect 360 1710 480 1755
rect 615 1740 690 1755
rect 750 1740 810 1755
rect 945 1740 1005 1755
rect 1080 1740 1155 1755
rect 1275 1740 1350 1755
rect 1410 1740 1485 1755
rect 1800 1740 2295 1770
rect 2370 1770 2490 1785
rect 2370 1755 2505 1770
rect 600 1725 675 1740
rect 765 1725 840 1740
rect 930 1725 990 1740
rect 1095 1725 1170 1740
rect 1260 1725 1335 1740
rect 1425 1725 1500 1740
rect 585 1710 660 1725
rect 780 1710 855 1725
rect 915 1710 975 1725
rect 1110 1710 1185 1725
rect 1245 1710 1320 1725
rect 1440 1710 1515 1725
rect 1785 1710 2295 1740
rect 2385 1725 2505 1755
rect 2385 1710 2520 1725
rect 345 1650 465 1710
rect 570 1695 645 1710
rect 795 1695 870 1710
rect 900 1695 960 1710
rect 1125 1695 1200 1710
rect 1230 1695 1305 1710
rect 1455 1695 1530 1710
rect 1800 1695 2295 1710
rect 555 1680 630 1695
rect 810 1680 945 1695
rect 1140 1680 1290 1695
rect 1470 1680 1545 1695
rect 1815 1680 2280 1695
rect 540 1665 600 1680
rect 825 1665 930 1680
rect 1155 1665 1275 1680
rect 1485 1665 1560 1680
rect 1830 1665 2280 1680
rect 2400 1665 2520 1710
rect 525 1650 585 1665
rect 330 1575 450 1650
rect 525 1635 600 1650
rect 840 1635 930 1665
rect 1170 1635 1260 1665
rect 1500 1635 1560 1665
rect 1740 1650 1755 1665
rect 1860 1650 2280 1665
rect 540 1620 600 1635
rect 825 1620 930 1635
rect 1155 1620 1275 1635
rect 1485 1620 1560 1635
rect 1725 1635 1770 1650
rect 1725 1620 1785 1635
rect 1875 1620 2280 1650
rect 555 1605 630 1620
rect 810 1605 945 1620
rect 1140 1605 1290 1620
rect 1470 1605 1545 1620
rect 1710 1605 1800 1620
rect 1890 1605 2010 1620
rect 2025 1605 2280 1620
rect 2415 1650 2520 1665
rect 570 1590 645 1605
rect 795 1590 870 1605
rect 900 1590 960 1605
rect 1125 1590 1200 1605
rect 1230 1590 1305 1605
rect 1455 1590 1530 1605
rect 1695 1590 1815 1605
rect 1905 1590 1965 1605
rect 2025 1590 2265 1605
rect 2415 1590 2535 1650
rect 585 1575 660 1590
rect 780 1575 855 1590
rect 915 1575 975 1590
rect 1110 1575 1185 1590
rect 1245 1575 1320 1590
rect 1440 1575 1515 1590
rect 1680 1575 1830 1590
rect 1920 1575 1935 1590
rect 2025 1575 2250 1590
rect 315 1560 435 1575
rect 600 1560 675 1575
rect 765 1560 840 1575
rect 930 1560 990 1575
rect 1095 1560 1170 1575
rect 1260 1560 1335 1575
rect 1425 1560 1500 1575
rect 1665 1560 1845 1575
rect 300 1530 435 1560
rect 615 1545 690 1560
rect 750 1545 810 1560
rect 945 1545 1005 1560
rect 1080 1545 1155 1560
rect 1275 1545 1350 1560
rect 1410 1545 1485 1560
rect 1650 1545 1860 1560
rect 2025 1545 2235 1575
rect 2430 1560 2535 1590
rect 630 1530 705 1545
rect 735 1530 795 1545
rect 960 1530 1035 1545
rect 1065 1530 1140 1545
rect 1290 1530 1365 1545
rect 1395 1530 1470 1545
rect 1620 1530 1845 1545
rect 2025 1530 2220 1545
rect 285 1515 435 1530
rect 645 1515 780 1530
rect 975 1515 1125 1530
rect 1305 1515 1455 1530
rect 1605 1515 1830 1530
rect 2025 1515 2205 1530
rect 270 1485 435 1515
rect 660 1500 765 1515
rect 990 1500 1110 1515
rect 1320 1500 1440 1515
rect 1590 1500 1815 1515
rect 2025 1500 2190 1515
rect 675 1485 750 1500
rect 255 1455 300 1485
rect 240 1425 285 1455
rect 225 1395 270 1425
rect 210 1380 255 1395
rect 195 1365 255 1380
rect 195 1335 240 1365
rect 180 1320 240 1335
rect 180 1290 225 1320
rect 315 1290 435 1485
rect 690 1470 765 1485
rect 1005 1470 1095 1500
rect 1335 1485 1425 1500
rect 1575 1485 1800 1500
rect 1335 1470 1410 1485
rect 1560 1470 1785 1485
rect 2025 1470 2175 1500
rect 705 1455 780 1470
rect 990 1455 1110 1470
rect 1320 1455 1395 1470
rect 1545 1455 1770 1470
rect 2025 1455 2160 1470
rect 720 1440 795 1455
rect 975 1440 1125 1455
rect 1305 1440 1380 1455
rect 1530 1440 1755 1455
rect 735 1425 795 1440
rect 960 1425 1035 1440
rect 1065 1425 1125 1440
rect 1290 1425 1365 1440
rect 1515 1425 1740 1440
rect 2025 1425 2145 1455
rect 750 1410 810 1425
rect 945 1410 1020 1425
rect 1080 1410 1140 1425
rect 1275 1410 1350 1425
rect 1500 1410 1725 1425
rect 2025 1410 2130 1425
rect 765 1395 840 1410
rect 930 1395 1005 1410
rect 1095 1395 1155 1410
rect 1260 1395 1335 1410
rect 1470 1395 1695 1410
rect 1785 1395 1815 1410
rect 2025 1395 2115 1410
rect 780 1380 855 1395
rect 915 1380 990 1395
rect 1110 1380 1170 1395
rect 1245 1380 1320 1395
rect 1455 1380 1680 1395
rect 1770 1380 1830 1395
rect 795 1365 870 1380
rect 900 1365 975 1380
rect 1125 1365 1185 1380
rect 1230 1365 1305 1380
rect 1440 1365 1665 1380
rect 1755 1365 1845 1380
rect 2025 1365 2100 1395
rect 810 1350 960 1365
rect 1140 1350 1290 1365
rect 1410 1350 1650 1365
rect 1740 1350 1860 1365
rect 2025 1350 2085 1365
rect 825 1335 945 1350
rect 1155 1335 1275 1350
rect 1395 1335 1620 1350
rect 1725 1335 1785 1350
rect 1800 1335 1875 1350
rect 2025 1335 2070 1350
rect 840 1320 930 1335
rect 1170 1320 1260 1335
rect 1380 1320 1605 1335
rect 1710 1320 1770 1335
rect 1815 1320 1890 1335
rect 2025 1320 2055 1335
rect 855 1305 915 1320
rect 1185 1305 1245 1320
rect 1350 1305 1590 1320
rect 1695 1305 1755 1320
rect 1830 1305 1905 1320
rect 2025 1305 2040 1320
rect 870 1290 885 1305
rect 1200 1290 1215 1305
rect 1335 1290 1560 1305
rect 1680 1290 1740 1305
rect 1860 1290 1920 1305
rect 165 1230 225 1290
rect 330 1260 435 1290
rect 1305 1275 1545 1290
rect 1665 1275 1725 1290
rect 1875 1275 1935 1290
rect 2430 1275 2550 1560
rect 1290 1260 1515 1275
rect 1650 1260 1710 1275
rect 1890 1260 1950 1275
rect 165 1170 210 1230
rect 330 1200 450 1260
rect 1260 1245 1500 1260
rect 1620 1245 1695 1260
rect 1905 1245 1965 1260
rect 2430 1245 2535 1275
rect 1245 1230 1470 1245
rect 1605 1230 1680 1245
rect 1215 1215 1455 1230
rect 1605 1215 1665 1230
rect 1200 1200 1440 1215
rect 1590 1200 1680 1215
rect 1920 1200 1980 1245
rect 345 1185 450 1200
rect 1170 1185 1410 1200
rect 1575 1185 1695 1200
rect 1905 1185 1965 1200
rect 2415 1185 2535 1245
rect 165 1110 225 1170
rect 345 1140 465 1185
rect 1155 1170 1380 1185
rect 1560 1170 1620 1185
rect 1635 1170 1710 1185
rect 1890 1170 1950 1185
rect 2415 1170 2520 1185
rect 1125 1155 1365 1170
rect 1545 1155 1605 1170
rect 1650 1155 1725 1170
rect 1875 1155 1935 1170
rect 1095 1140 1335 1155
rect 1530 1140 1590 1155
rect 1665 1140 1740 1155
rect 1860 1140 1920 1155
rect 360 1125 465 1140
rect 1080 1125 1305 1140
rect 1515 1125 1575 1140
rect 1680 1125 1755 1140
rect 1830 1125 1905 1140
rect 2400 1125 2520 1170
rect 165 1095 240 1110
rect 180 1080 240 1095
rect 360 1080 480 1125
rect 1050 1110 1275 1125
rect 1500 1110 1560 1125
rect 1695 1110 1770 1125
rect 1815 1110 1890 1125
rect 1020 1095 1260 1110
rect 1485 1095 1545 1110
rect 1710 1095 1785 1110
rect 1800 1095 1875 1110
rect 990 1080 1230 1095
rect 1470 1080 1530 1095
rect 1725 1080 1860 1095
rect 2385 1080 2505 1125
rect 180 1065 255 1080
rect 180 1050 270 1065
rect 195 1035 270 1050
rect 375 1050 495 1080
rect 960 1065 1200 1080
rect 1455 1065 1515 1080
rect 1740 1065 1845 1080
rect 930 1050 1170 1065
rect 1440 1050 1500 1065
rect 1755 1050 1830 1065
rect 375 1035 510 1050
rect 900 1035 1140 1050
rect 1440 1035 1515 1050
rect 1740 1035 1845 1050
rect 2370 1035 2490 1080
rect 210 1020 300 1035
rect 420 1020 510 1035
rect 855 1020 1110 1035
rect 1455 1020 1530 1035
rect 1725 1020 1860 1035
rect 210 1005 315 1020
rect 480 1005 510 1020
rect 825 1005 1080 1020
rect 1470 1005 1545 1020
rect 1725 1005 1785 1020
rect 1800 1005 1875 1020
rect 2355 1005 2475 1035
rect 225 990 330 1005
rect 780 990 1050 1005
rect 1485 990 1560 1005
rect 1710 990 1770 1005
rect 1815 990 1890 1005
rect 2340 990 2475 1005
rect 240 975 360 990
rect 735 975 1020 990
rect 1500 975 1575 990
rect 1695 975 1755 990
rect 1830 975 1905 990
rect 2340 975 2460 990
rect 255 960 405 975
rect 690 960 975 975
rect 1515 960 1590 975
rect 1680 960 1740 975
rect 1845 960 1920 975
rect 2325 960 2460 975
rect 285 945 480 960
rect 600 945 945 960
rect 1530 945 1605 960
rect 1665 945 1725 960
rect 1860 945 1935 960
rect 2325 945 2445 960
rect 300 930 900 945
rect 1545 930 1620 945
rect 1650 930 1710 945
rect 1875 930 1950 945
rect 2310 930 2445 945
rect 330 915 855 930
rect 1560 915 1695 930
rect 1890 915 1965 930
rect 2310 915 2430 930
rect 360 900 810 915
rect 1575 900 1680 915
rect 1905 900 1980 915
rect 390 885 750 900
rect 1590 885 1665 900
rect 465 870 675 885
rect 1590 870 1680 885
rect 1920 870 1980 900
rect 2295 900 2430 915
rect 2295 885 2415 900
rect 2280 870 2415 885
rect 1575 855 1695 870
rect 1905 855 1965 870
rect 1560 840 1620 855
rect 1635 840 1710 855
rect 1890 840 1950 855
rect 2265 840 2400 870
rect 2640 855 2655 870
rect 2625 840 2655 855
rect 1545 825 1605 840
rect 1650 825 1725 840
rect 1875 825 1935 840
rect 2250 825 2385 840
rect 1530 810 1590 825
rect 1665 810 1740 825
rect 1860 810 1920 825
rect 2235 810 2370 825
rect 2625 810 2670 840
rect 495 795 645 810
rect 1515 795 1575 810
rect 1680 795 1755 810
rect 1845 795 1905 810
rect 2220 795 2370 810
rect 2610 795 2685 810
rect 510 780 660 795
rect 1500 780 1560 795
rect 1695 780 1770 795
rect 1830 780 1890 795
rect 2220 780 2355 795
rect 2595 780 2700 795
rect 525 765 660 780
rect 1485 765 1545 780
rect 1710 765 1785 780
rect 1815 765 1875 780
rect 2205 765 2340 780
rect 2580 765 2715 780
rect 525 750 675 765
rect 1470 750 1530 765
rect 1725 750 1860 765
rect 2190 750 2340 765
rect 2550 750 2745 765
rect 540 735 690 750
rect 1455 735 1515 750
rect 1740 735 1845 750
rect 2175 735 2325 750
rect 2520 735 2775 750
rect 555 720 705 735
rect 1440 720 1500 735
rect 1755 720 1830 735
rect 2160 720 2310 735
rect 2565 720 2730 735
rect 570 705 720 720
rect 1440 705 1515 720
rect 1755 705 1815 720
rect 2145 705 2295 720
rect 2580 705 2700 720
rect 585 690 735 705
rect 1455 690 1530 705
rect 1740 690 1800 705
rect 2130 690 2295 705
rect 2595 690 2685 705
rect 600 675 750 690
rect 1470 675 1545 690
rect 1725 675 1785 690
rect 2115 675 2280 690
rect 2610 675 2670 690
rect 600 660 765 675
rect 1485 660 1560 675
rect 1710 660 1770 675
rect 2100 660 2265 675
rect 2625 660 2670 675
rect 630 645 780 660
rect 1500 645 1575 660
rect 1695 645 1755 660
rect 2085 645 2250 660
rect 2625 645 2655 660
rect 645 630 810 645
rect 1515 630 1590 645
rect 1680 630 1740 645
rect 2070 630 2235 645
rect 2640 630 2655 645
rect 660 615 825 630
rect 1530 615 1605 630
rect 1665 615 1725 630
rect 2040 615 2220 630
rect 660 600 840 615
rect 1545 600 1605 615
rect 1650 600 1710 615
rect 2025 600 2205 615
rect 675 585 870 600
rect 1560 585 1695 600
rect 2010 585 2190 600
rect 705 570 885 585
rect 1575 570 1680 585
rect 1980 570 2175 585
rect 720 555 915 570
rect 1590 555 1665 570
rect 1965 555 2145 570
rect 735 540 930 555
rect 1605 540 1650 555
rect 1935 540 2130 555
rect 750 525 960 540
rect 1905 525 2115 540
rect 780 510 990 525
rect 1875 510 2100 525
rect 795 495 1020 510
rect 1845 495 2070 510
rect 810 480 1065 495
rect 1800 480 2055 495
rect 840 465 1095 480
rect 1770 465 2025 480
rect 870 450 1155 465
rect 1725 450 1995 465
rect 900 435 1200 450
rect 1665 435 1980 450
rect 915 420 1290 435
rect 1575 420 1950 435
rect 945 405 1920 420
rect 975 390 1890 405
rect 1005 375 1860 390
rect 1050 360 1815 375
rect 1095 345 1770 360
rect 1155 330 1710 345
rect 1215 315 1650 330
rect 1320 300 1545 315
<< metal4 >>
rect 2775 2610 2850 2625
rect 2715 2595 2850 2610
rect 2670 2580 2835 2595
rect 2625 2565 2835 2580
rect 2580 2550 2835 2565
rect 2550 2535 2835 2550
rect 1275 2520 1590 2535
rect 2520 2520 2820 2535
rect 1185 2505 1680 2520
rect 2490 2505 2820 2520
rect 1125 2490 1740 2505
rect 2460 2490 2820 2505
rect 1080 2475 1785 2490
rect 2445 2475 2820 2490
rect 1035 2460 1830 2475
rect 2415 2460 2805 2475
rect 1005 2445 1860 2460
rect 2400 2445 2805 2460
rect 975 2430 1890 2445
rect 2370 2430 2805 2445
rect 240 2370 255 2430
rect 945 2415 1395 2430
rect 1470 2415 1920 2430
rect 2355 2415 2790 2430
rect 915 2400 1260 2415
rect 1605 2400 1950 2415
rect 2340 2400 2790 2415
rect 885 2385 1185 2400
rect 1680 2385 1980 2400
rect 2310 2385 2775 2400
rect 855 2370 1125 2385
rect 1740 2370 2010 2385
rect 2295 2370 2775 2385
rect 225 2340 270 2370
rect 840 2355 1080 2370
rect 1785 2355 2040 2370
rect 2280 2355 2775 2370
rect 810 2340 1050 2355
rect 1815 2340 2055 2355
rect 2265 2340 2430 2355
rect 2535 2340 2760 2355
rect 210 2325 285 2340
rect 780 2325 1005 2340
rect 1860 2325 2085 2340
rect 2235 2325 2415 2340
rect 2550 2325 2760 2340
rect 195 2310 285 2325
rect 765 2310 975 2325
rect 1890 2310 2100 2325
rect 2220 2310 2400 2325
rect 180 2295 300 2310
rect 750 2295 945 2310
rect 1920 2295 2115 2310
rect 2205 2295 2400 2310
rect 2565 2295 2745 2325
rect 180 2280 315 2295
rect 720 2280 930 2295
rect 1935 2280 2100 2295
rect 2190 2280 2400 2295
rect 150 2265 330 2280
rect 705 2265 900 2280
rect 1965 2265 2085 2280
rect 2175 2265 2400 2280
rect 2580 2280 2730 2295
rect 2580 2265 2715 2280
rect 135 2250 360 2265
rect 690 2250 870 2265
rect 1995 2250 2070 2265
rect 2160 2250 2400 2265
rect 120 2235 375 2250
rect 675 2235 855 2250
rect 2010 2235 2070 2250
rect 2145 2235 2400 2250
rect 90 2220 405 2235
rect 660 2220 840 2235
rect 2025 2220 2055 2235
rect 2130 2220 2400 2235
rect 2565 2250 2715 2265
rect 2565 2220 2700 2250
rect 15 2205 465 2220
rect 645 2205 810 2220
rect 2115 2205 2415 2220
rect 2550 2205 2685 2220
rect 90 2190 405 2205
rect 630 2190 795 2205
rect 2100 2190 2430 2205
rect 2535 2190 2670 2205
rect 120 2175 375 2190
rect 615 2175 780 2190
rect 2100 2175 2475 2190
rect 2505 2175 2670 2190
rect 135 2160 345 2175
rect 600 2160 765 2175
rect 2085 2160 2655 2175
rect 165 2145 330 2160
rect 585 2145 750 2160
rect 2070 2145 2640 2160
rect 180 2130 315 2145
rect 570 2130 735 2145
rect 2055 2130 2625 2145
rect 195 2115 300 2130
rect 570 2115 720 2130
rect 2040 2115 2625 2130
rect 195 2100 285 2115
rect 555 2100 705 2115
rect 2025 2100 2610 2115
rect 210 2085 285 2100
rect 540 2085 690 2100
rect 1995 2085 2595 2100
rect 225 2055 270 2085
rect 525 2070 675 2085
rect 1845 2070 2580 2085
rect 525 2055 660 2070
rect 1800 2055 2565 2070
rect 240 1995 255 2055
rect 510 2040 645 2055
rect 1785 2040 2565 2055
rect 495 2025 645 2040
rect 1770 2025 2550 2040
rect 495 2010 630 2025
rect 1755 2010 2535 2025
rect 480 1995 615 2010
rect 1725 1995 2520 2010
rect 465 1965 600 1995
rect 1710 1980 2505 1995
rect 1695 1965 2490 1980
rect 450 1950 585 1965
rect 1665 1950 2475 1965
rect 450 1935 570 1950
rect 1650 1935 2460 1950
rect 435 1920 570 1935
rect 1620 1920 2445 1935
rect 435 1905 555 1920
rect 1605 1905 2430 1920
rect 420 1890 555 1905
rect 1590 1890 2415 1905
rect 420 1875 540 1890
rect 1575 1875 2385 1890
rect 405 1860 540 1875
rect 1545 1860 2370 1875
rect 405 1845 525 1860
rect 1530 1845 2355 1860
rect 2445 1845 2460 1860
rect 390 1830 525 1845
rect 1515 1830 2340 1845
rect 2430 1830 2475 1845
rect 390 1800 510 1830
rect 690 1815 735 1830
rect 1020 1815 1080 1830
rect 1350 1815 1410 1830
rect 1665 1815 2325 1830
rect 2415 1815 2475 1830
rect 675 1800 750 1815
rect 1005 1800 1095 1815
rect 1335 1800 1425 1815
rect 375 1755 495 1800
rect 660 1785 765 1800
rect 990 1785 1110 1800
rect 1320 1785 1440 1800
rect 645 1770 780 1785
rect 975 1770 1125 1785
rect 1305 1770 1455 1785
rect 1815 1770 2295 1815
rect 2400 1800 2490 1815
rect 2385 1785 2490 1800
rect 630 1755 705 1770
rect 735 1755 795 1770
rect 960 1755 1035 1770
rect 1065 1755 1140 1770
rect 1290 1755 1365 1770
rect 1395 1755 1470 1770
rect 360 1710 480 1755
rect 615 1740 690 1755
rect 750 1740 810 1755
rect 945 1740 1005 1755
rect 1080 1740 1155 1755
rect 1275 1740 1350 1755
rect 1410 1740 1485 1755
rect 1800 1740 2295 1770
rect 2370 1770 2490 1785
rect 2370 1755 2505 1770
rect 600 1725 675 1740
rect 765 1725 840 1740
rect 930 1725 990 1740
rect 1095 1725 1170 1740
rect 1260 1725 1335 1740
rect 1425 1725 1500 1740
rect 585 1710 660 1725
rect 780 1710 855 1725
rect 915 1710 975 1725
rect 1110 1710 1185 1725
rect 1245 1710 1320 1725
rect 1440 1710 1515 1725
rect 1785 1710 2295 1740
rect 2385 1725 2505 1755
rect 2385 1710 2520 1725
rect 345 1650 465 1710
rect 570 1695 645 1710
rect 795 1695 870 1710
rect 900 1695 960 1710
rect 1125 1695 1200 1710
rect 1230 1695 1305 1710
rect 1455 1695 1530 1710
rect 1800 1695 2295 1710
rect 555 1680 630 1695
rect 810 1680 945 1695
rect 1140 1680 1290 1695
rect 1470 1680 1545 1695
rect 1815 1680 2280 1695
rect 540 1665 600 1680
rect 825 1665 930 1680
rect 1155 1665 1275 1680
rect 1485 1665 1560 1680
rect 1830 1665 2280 1680
rect 2400 1665 2520 1710
rect 525 1650 585 1665
rect 330 1575 450 1650
rect 525 1635 600 1650
rect 840 1635 930 1665
rect 1170 1635 1260 1665
rect 1500 1635 1560 1665
rect 1740 1650 1755 1665
rect 1860 1650 2280 1665
rect 540 1620 600 1635
rect 825 1620 930 1635
rect 1155 1620 1275 1635
rect 1485 1620 1560 1635
rect 1725 1635 1770 1650
rect 1725 1620 1785 1635
rect 1875 1620 2280 1650
rect 555 1605 630 1620
rect 810 1605 945 1620
rect 1140 1605 1290 1620
rect 1470 1605 1545 1620
rect 1710 1605 1800 1620
rect 1890 1605 2010 1620
rect 2025 1605 2280 1620
rect 2415 1650 2520 1665
rect 570 1590 645 1605
rect 795 1590 870 1605
rect 900 1590 960 1605
rect 1125 1590 1200 1605
rect 1230 1590 1305 1605
rect 1455 1590 1530 1605
rect 1695 1590 1815 1605
rect 1905 1590 1965 1605
rect 2025 1590 2265 1605
rect 2415 1590 2535 1650
rect 585 1575 660 1590
rect 780 1575 855 1590
rect 915 1575 975 1590
rect 1110 1575 1185 1590
rect 1245 1575 1320 1590
rect 1440 1575 1515 1590
rect 1680 1575 1830 1590
rect 1920 1575 1935 1590
rect 2025 1575 2250 1590
rect 315 1560 435 1575
rect 600 1560 675 1575
rect 765 1560 840 1575
rect 930 1560 990 1575
rect 1095 1560 1170 1575
rect 1260 1560 1335 1575
rect 1425 1560 1500 1575
rect 1665 1560 1845 1575
rect 300 1530 435 1560
rect 615 1545 690 1560
rect 750 1545 810 1560
rect 945 1545 1005 1560
rect 1080 1545 1155 1560
rect 1275 1545 1350 1560
rect 1410 1545 1485 1560
rect 1650 1545 1860 1560
rect 2025 1545 2235 1575
rect 2430 1560 2535 1590
rect 630 1530 705 1545
rect 735 1530 795 1545
rect 960 1530 1035 1545
rect 1065 1530 1140 1545
rect 1290 1530 1365 1545
rect 1395 1530 1470 1545
rect 1620 1530 1845 1545
rect 2025 1530 2220 1545
rect 285 1515 435 1530
rect 645 1515 780 1530
rect 975 1515 1125 1530
rect 1305 1515 1455 1530
rect 1605 1515 1830 1530
rect 2025 1515 2205 1530
rect 270 1485 435 1515
rect 660 1500 765 1515
rect 990 1500 1110 1515
rect 1320 1500 1440 1515
rect 1590 1500 1815 1515
rect 2025 1500 2190 1515
rect 675 1485 750 1500
rect 255 1455 300 1485
rect 240 1425 285 1455
rect 225 1395 270 1425
rect 210 1380 255 1395
rect 195 1365 255 1380
rect 195 1335 240 1365
rect 180 1320 240 1335
rect 180 1290 225 1320
rect 315 1290 435 1485
rect 690 1470 765 1485
rect 1005 1470 1095 1500
rect 1335 1485 1425 1500
rect 1575 1485 1800 1500
rect 1335 1470 1410 1485
rect 1560 1470 1785 1485
rect 2025 1470 2175 1500
rect 705 1455 780 1470
rect 990 1455 1110 1470
rect 1320 1455 1395 1470
rect 1545 1455 1770 1470
rect 2025 1455 2160 1470
rect 720 1440 795 1455
rect 975 1440 1125 1455
rect 1305 1440 1380 1455
rect 1530 1440 1755 1455
rect 735 1425 795 1440
rect 960 1425 1035 1440
rect 1065 1425 1125 1440
rect 1290 1425 1365 1440
rect 1515 1425 1740 1440
rect 2025 1425 2145 1455
rect 750 1410 810 1425
rect 945 1410 1020 1425
rect 1080 1410 1140 1425
rect 1275 1410 1350 1425
rect 1500 1410 1725 1425
rect 2025 1410 2130 1425
rect 765 1395 840 1410
rect 930 1395 1005 1410
rect 1095 1395 1155 1410
rect 1260 1395 1335 1410
rect 1470 1395 1695 1410
rect 1785 1395 1815 1410
rect 2025 1395 2115 1410
rect 780 1380 855 1395
rect 915 1380 990 1395
rect 1110 1380 1170 1395
rect 1245 1380 1320 1395
rect 1455 1380 1680 1395
rect 1770 1380 1830 1395
rect 795 1365 870 1380
rect 900 1365 975 1380
rect 1125 1365 1185 1380
rect 1230 1365 1305 1380
rect 1440 1365 1665 1380
rect 1755 1365 1845 1380
rect 2025 1365 2100 1395
rect 810 1350 960 1365
rect 1140 1350 1290 1365
rect 1410 1350 1650 1365
rect 1740 1350 1860 1365
rect 2025 1350 2085 1365
rect 825 1335 945 1350
rect 1155 1335 1275 1350
rect 1395 1335 1620 1350
rect 1725 1335 1785 1350
rect 1800 1335 1875 1350
rect 2025 1335 2070 1350
rect 840 1320 930 1335
rect 1170 1320 1260 1335
rect 1380 1320 1605 1335
rect 1710 1320 1770 1335
rect 1815 1320 1890 1335
rect 2025 1320 2055 1335
rect 855 1305 915 1320
rect 1185 1305 1245 1320
rect 1350 1305 1590 1320
rect 1695 1305 1755 1320
rect 1830 1305 1905 1320
rect 2025 1305 2040 1320
rect 870 1290 885 1305
rect 1200 1290 1215 1305
rect 1335 1290 1560 1305
rect 1680 1290 1740 1305
rect 1860 1290 1920 1305
rect 165 1230 225 1290
rect 330 1260 435 1290
rect 1305 1275 1545 1290
rect 1665 1275 1725 1290
rect 1875 1275 1935 1290
rect 2430 1275 2550 1560
rect 1290 1260 1515 1275
rect 1650 1260 1710 1275
rect 1890 1260 1950 1275
rect 165 1170 210 1230
rect 330 1200 450 1260
rect 1260 1245 1500 1260
rect 1620 1245 1695 1260
rect 1905 1245 1965 1260
rect 2430 1245 2535 1275
rect 1245 1230 1470 1245
rect 1605 1230 1680 1245
rect 1215 1215 1455 1230
rect 1605 1215 1665 1230
rect 1200 1200 1440 1215
rect 1590 1200 1680 1215
rect 1920 1200 1980 1245
rect 345 1185 450 1200
rect 1170 1185 1410 1200
rect 1575 1185 1695 1200
rect 1905 1185 1965 1200
rect 2415 1185 2535 1245
rect 165 1110 225 1170
rect 345 1140 465 1185
rect 1155 1170 1380 1185
rect 1560 1170 1620 1185
rect 1635 1170 1710 1185
rect 1890 1170 1950 1185
rect 2415 1170 2520 1185
rect 1125 1155 1365 1170
rect 1545 1155 1605 1170
rect 1650 1155 1725 1170
rect 1875 1155 1935 1170
rect 1095 1140 1335 1155
rect 1530 1140 1590 1155
rect 1665 1140 1740 1155
rect 1860 1140 1920 1155
rect 360 1125 465 1140
rect 1080 1125 1305 1140
rect 1515 1125 1575 1140
rect 1680 1125 1755 1140
rect 1830 1125 1905 1140
rect 2400 1125 2520 1170
rect 165 1095 240 1110
rect 180 1080 240 1095
rect 360 1080 480 1125
rect 1050 1110 1275 1125
rect 1500 1110 1560 1125
rect 1695 1110 1770 1125
rect 1815 1110 1890 1125
rect 1020 1095 1260 1110
rect 1485 1095 1545 1110
rect 1710 1095 1785 1110
rect 1800 1095 1875 1110
rect 990 1080 1230 1095
rect 1470 1080 1530 1095
rect 1725 1080 1860 1095
rect 2385 1080 2505 1125
rect 180 1065 255 1080
rect 180 1050 270 1065
rect 195 1035 270 1050
rect 375 1050 495 1080
rect 960 1065 1200 1080
rect 1455 1065 1515 1080
rect 1740 1065 1845 1080
rect 930 1050 1170 1065
rect 1440 1050 1500 1065
rect 1755 1050 1830 1065
rect 375 1035 510 1050
rect 900 1035 1140 1050
rect 1440 1035 1515 1050
rect 1740 1035 1845 1050
rect 2370 1035 2490 1080
rect 210 1020 300 1035
rect 420 1020 510 1035
rect 855 1020 1110 1035
rect 1455 1020 1530 1035
rect 1725 1020 1860 1035
rect 210 1005 315 1020
rect 480 1005 510 1020
rect 825 1005 1080 1020
rect 1470 1005 1545 1020
rect 1725 1005 1785 1020
rect 1800 1005 1875 1020
rect 2355 1005 2475 1035
rect 225 990 330 1005
rect 780 990 1050 1005
rect 1485 990 1560 1005
rect 1710 990 1770 1005
rect 1815 990 1890 1005
rect 2340 990 2475 1005
rect 240 975 360 990
rect 735 975 1020 990
rect 1500 975 1575 990
rect 1695 975 1755 990
rect 1830 975 1905 990
rect 2340 975 2460 990
rect 255 960 405 975
rect 690 960 975 975
rect 1515 960 1590 975
rect 1680 960 1740 975
rect 1845 960 1920 975
rect 2325 960 2460 975
rect 285 945 480 960
rect 600 945 945 960
rect 1530 945 1605 960
rect 1665 945 1725 960
rect 1860 945 1935 960
rect 2325 945 2445 960
rect 300 930 900 945
rect 1545 930 1620 945
rect 1650 930 1710 945
rect 1875 930 1950 945
rect 2310 930 2445 945
rect 330 915 855 930
rect 1560 915 1695 930
rect 1890 915 1965 930
rect 2310 915 2430 930
rect 360 900 810 915
rect 1575 900 1680 915
rect 1905 900 1980 915
rect 390 885 750 900
rect 1590 885 1665 900
rect 465 870 675 885
rect 1590 870 1680 885
rect 1920 870 1980 900
rect 2295 900 2430 915
rect 2295 885 2415 900
rect 2280 870 2415 885
rect 1575 855 1695 870
rect 1905 855 1965 870
rect 1560 840 1620 855
rect 1635 840 1710 855
rect 1890 840 1950 855
rect 2265 840 2400 870
rect 2640 855 2655 870
rect 2625 840 2655 855
rect 1545 825 1605 840
rect 1650 825 1725 840
rect 1875 825 1935 840
rect 2250 825 2385 840
rect 1530 810 1590 825
rect 1665 810 1740 825
rect 1860 810 1920 825
rect 2235 810 2370 825
rect 2625 810 2670 840
rect 495 795 645 810
rect 1515 795 1575 810
rect 1680 795 1755 810
rect 1845 795 1905 810
rect 2220 795 2370 810
rect 2610 795 2685 810
rect 510 780 660 795
rect 1500 780 1560 795
rect 1695 780 1770 795
rect 1830 780 1890 795
rect 2220 780 2355 795
rect 2595 780 2700 795
rect 525 765 660 780
rect 1485 765 1545 780
rect 1710 765 1785 780
rect 1815 765 1875 780
rect 2205 765 2340 780
rect 2580 765 2715 780
rect 525 750 675 765
rect 1470 750 1530 765
rect 1725 750 1860 765
rect 2190 750 2340 765
rect 2550 750 2745 765
rect 540 735 690 750
rect 1455 735 1515 750
rect 1740 735 1845 750
rect 2175 735 2325 750
rect 2520 735 2775 750
rect 555 720 705 735
rect 1440 720 1500 735
rect 1755 720 1830 735
rect 2160 720 2310 735
rect 2565 720 2730 735
rect 570 705 720 720
rect 1440 705 1515 720
rect 1755 705 1815 720
rect 2145 705 2295 720
rect 2580 705 2700 720
rect 585 690 735 705
rect 1455 690 1530 705
rect 1740 690 1800 705
rect 2130 690 2295 705
rect 2595 690 2685 705
rect 600 675 750 690
rect 1470 675 1545 690
rect 1725 675 1785 690
rect 2115 675 2280 690
rect 2610 675 2670 690
rect 600 660 765 675
rect 1485 660 1560 675
rect 1710 660 1770 675
rect 2100 660 2265 675
rect 2625 660 2670 675
rect 630 645 780 660
rect 1500 645 1575 660
rect 1695 645 1755 660
rect 2085 645 2250 660
rect 2625 645 2655 660
rect 645 630 810 645
rect 1515 630 1590 645
rect 1680 630 1740 645
rect 2070 630 2235 645
rect 2640 630 2655 645
rect 660 615 825 630
rect 1530 615 1605 630
rect 1665 615 1725 630
rect 2040 615 2220 630
rect 660 600 840 615
rect 1545 600 1605 615
rect 1650 600 1710 615
rect 2025 600 2205 615
rect 675 585 870 600
rect 1560 585 1695 600
rect 2010 585 2190 600
rect 705 570 885 585
rect 1575 570 1680 585
rect 1980 570 2175 585
rect 720 555 915 570
rect 1590 555 1665 570
rect 1965 555 2145 570
rect 735 540 930 555
rect 1605 540 1650 555
rect 1935 540 2130 555
rect 750 525 960 540
rect 1905 525 2115 540
rect 780 510 990 525
rect 1875 510 2100 525
rect 795 495 1020 510
rect 1845 495 2070 510
rect 810 480 1065 495
rect 1800 480 2055 495
rect 840 465 1095 480
rect 1770 465 2025 480
rect 870 450 1155 465
rect 1725 450 1995 465
rect 900 435 1200 450
rect 1665 435 1980 450
rect 915 420 1290 435
rect 1575 420 1950 435
rect 945 405 1920 420
rect 975 390 1890 405
rect 1005 375 1860 390
rect 1050 360 1815 375
rect 1095 345 1770 360
rect 1155 330 1710 345
rect 1215 315 1650 330
rect 1320 300 1545 315
<< metal5 >>
rect 2775 2610 2850 2625
rect 2715 2595 2850 2610
rect 2670 2580 2835 2595
rect 2625 2565 2835 2580
rect 2580 2550 2835 2565
rect 2550 2535 2835 2550
rect 1275 2520 1590 2535
rect 2520 2520 2820 2535
rect 1185 2505 1680 2520
rect 2490 2505 2820 2520
rect 1125 2490 1740 2505
rect 2460 2490 2820 2505
rect 1080 2475 1785 2490
rect 2445 2475 2820 2490
rect 1035 2460 1830 2475
rect 2415 2460 2805 2475
rect 1005 2445 1860 2460
rect 2400 2445 2805 2460
rect 975 2430 1890 2445
rect 2370 2430 2805 2445
rect 240 2370 255 2430
rect 945 2415 1395 2430
rect 1470 2415 1920 2430
rect 2355 2415 2790 2430
rect 915 2400 1260 2415
rect 1605 2400 1950 2415
rect 2340 2400 2790 2415
rect 885 2385 1185 2400
rect 1680 2385 1980 2400
rect 2310 2385 2775 2400
rect 855 2370 1125 2385
rect 1740 2370 2010 2385
rect 2295 2370 2775 2385
rect 225 2340 270 2370
rect 840 2355 1080 2370
rect 1785 2355 2040 2370
rect 2280 2355 2775 2370
rect 810 2340 1050 2355
rect 1815 2340 2055 2355
rect 2265 2340 2430 2355
rect 2535 2340 2760 2355
rect 210 2325 285 2340
rect 780 2325 1005 2340
rect 1860 2325 2085 2340
rect 2235 2325 2415 2340
rect 2550 2325 2760 2340
rect 195 2310 285 2325
rect 765 2310 975 2325
rect 1890 2310 2100 2325
rect 2220 2310 2400 2325
rect 180 2295 300 2310
rect 750 2295 945 2310
rect 1920 2295 2115 2310
rect 2205 2295 2400 2310
rect 2565 2295 2745 2325
rect 180 2280 315 2295
rect 720 2280 930 2295
rect 1935 2280 2100 2295
rect 2190 2280 2400 2295
rect 150 2265 330 2280
rect 705 2265 900 2280
rect 1965 2265 2085 2280
rect 2175 2265 2400 2280
rect 2580 2280 2730 2295
rect 2580 2265 2715 2280
rect 135 2250 360 2265
rect 690 2250 870 2265
rect 1995 2250 2070 2265
rect 2160 2250 2400 2265
rect 120 2235 375 2250
rect 675 2235 855 2250
rect 2010 2235 2070 2250
rect 2145 2235 2400 2250
rect 90 2220 405 2235
rect 660 2220 840 2235
rect 2025 2220 2055 2235
rect 2130 2220 2400 2235
rect 2565 2250 2715 2265
rect 2565 2220 2700 2250
rect 15 2205 465 2220
rect 645 2205 810 2220
rect 2115 2205 2415 2220
rect 2550 2205 2685 2220
rect 90 2190 405 2205
rect 630 2190 795 2205
rect 2100 2190 2430 2205
rect 2535 2190 2670 2205
rect 120 2175 375 2190
rect 615 2175 780 2190
rect 2100 2175 2475 2190
rect 2505 2175 2670 2190
rect 135 2160 345 2175
rect 600 2160 765 2175
rect 2085 2160 2655 2175
rect 165 2145 330 2160
rect 585 2145 750 2160
rect 2070 2145 2640 2160
rect 180 2130 315 2145
rect 570 2130 735 2145
rect 2055 2130 2625 2145
rect 195 2115 300 2130
rect 570 2115 720 2130
rect 2040 2115 2625 2130
rect 195 2100 285 2115
rect 555 2100 705 2115
rect 2025 2100 2610 2115
rect 210 2085 285 2100
rect 540 2085 690 2100
rect 1995 2085 2595 2100
rect 225 2055 270 2085
rect 525 2070 675 2085
rect 1845 2070 2580 2085
rect 525 2055 660 2070
rect 1800 2055 2565 2070
rect 240 1995 255 2055
rect 510 2040 645 2055
rect 1785 2040 2565 2055
rect 495 2025 645 2040
rect 1770 2025 2550 2040
rect 495 2010 630 2025
rect 1755 2010 2535 2025
rect 480 1995 615 2010
rect 1725 1995 2520 2010
rect 465 1965 600 1995
rect 1710 1980 2505 1995
rect 1695 1965 2490 1980
rect 450 1950 585 1965
rect 1665 1950 2475 1965
rect 450 1935 570 1950
rect 1650 1935 2460 1950
rect 435 1920 570 1935
rect 1620 1920 2445 1935
rect 435 1905 555 1920
rect 1605 1905 2430 1920
rect 420 1890 555 1905
rect 1590 1890 2415 1905
rect 420 1875 540 1890
rect 1575 1875 2385 1890
rect 405 1860 540 1875
rect 1545 1860 2370 1875
rect 405 1845 525 1860
rect 1530 1845 2355 1860
rect 2445 1845 2460 1860
rect 390 1830 525 1845
rect 1515 1830 2340 1845
rect 2430 1830 2475 1845
rect 390 1800 510 1830
rect 690 1815 735 1830
rect 1020 1815 1080 1830
rect 1350 1815 1410 1830
rect 1665 1815 2325 1830
rect 2415 1815 2475 1830
rect 675 1800 750 1815
rect 1005 1800 1095 1815
rect 1335 1800 1425 1815
rect 375 1755 495 1800
rect 660 1785 765 1800
rect 990 1785 1110 1800
rect 1320 1785 1440 1800
rect 645 1770 780 1785
rect 975 1770 1125 1785
rect 1305 1770 1455 1785
rect 1815 1770 2295 1815
rect 2400 1800 2490 1815
rect 2385 1785 2490 1800
rect 630 1755 705 1770
rect 735 1755 795 1770
rect 960 1755 1035 1770
rect 1065 1755 1140 1770
rect 1290 1755 1365 1770
rect 1395 1755 1470 1770
rect 360 1710 480 1755
rect 615 1740 690 1755
rect 750 1740 810 1755
rect 945 1740 1005 1755
rect 1080 1740 1155 1755
rect 1275 1740 1350 1755
rect 1410 1740 1485 1755
rect 1800 1740 2295 1770
rect 2370 1770 2490 1785
rect 2370 1755 2505 1770
rect 600 1725 675 1740
rect 765 1725 840 1740
rect 930 1725 990 1740
rect 1095 1725 1170 1740
rect 1260 1725 1335 1740
rect 1425 1725 1500 1740
rect 585 1710 660 1725
rect 780 1710 855 1725
rect 915 1710 975 1725
rect 1110 1710 1185 1725
rect 1245 1710 1320 1725
rect 1440 1710 1515 1725
rect 1785 1710 2295 1740
rect 2385 1725 2505 1755
rect 2385 1710 2520 1725
rect 345 1650 465 1710
rect 570 1695 645 1710
rect 795 1695 870 1710
rect 900 1695 960 1710
rect 1125 1695 1200 1710
rect 1230 1695 1305 1710
rect 1455 1695 1530 1710
rect 1800 1695 2295 1710
rect 555 1680 630 1695
rect 810 1680 945 1695
rect 1140 1680 1290 1695
rect 1470 1680 1545 1695
rect 1815 1680 2280 1695
rect 540 1665 600 1680
rect 825 1665 930 1680
rect 1155 1665 1275 1680
rect 1485 1665 1560 1680
rect 1830 1665 2280 1680
rect 2400 1665 2520 1710
rect 525 1650 585 1665
rect 330 1575 450 1650
rect 525 1635 600 1650
rect 840 1635 930 1665
rect 1170 1635 1260 1665
rect 1500 1635 1560 1665
rect 1740 1650 1755 1665
rect 1860 1650 2280 1665
rect 540 1620 600 1635
rect 825 1620 930 1635
rect 1155 1620 1275 1635
rect 1485 1620 1560 1635
rect 1725 1635 1770 1650
rect 1725 1620 1785 1635
rect 1875 1620 2280 1650
rect 555 1605 630 1620
rect 810 1605 945 1620
rect 1140 1605 1290 1620
rect 1470 1605 1545 1620
rect 1710 1605 1800 1620
rect 1890 1605 2010 1620
rect 2025 1605 2280 1620
rect 2415 1650 2520 1665
rect 570 1590 645 1605
rect 795 1590 870 1605
rect 900 1590 960 1605
rect 1125 1590 1200 1605
rect 1230 1590 1305 1605
rect 1455 1590 1530 1605
rect 1695 1590 1815 1605
rect 1905 1590 1965 1605
rect 2025 1590 2265 1605
rect 2415 1590 2535 1650
rect 585 1575 660 1590
rect 780 1575 855 1590
rect 915 1575 975 1590
rect 1110 1575 1185 1590
rect 1245 1575 1320 1590
rect 1440 1575 1515 1590
rect 1680 1575 1830 1590
rect 1920 1575 1935 1590
rect 2025 1575 2250 1590
rect 315 1560 435 1575
rect 600 1560 675 1575
rect 765 1560 840 1575
rect 930 1560 990 1575
rect 1095 1560 1170 1575
rect 1260 1560 1335 1575
rect 1425 1560 1500 1575
rect 1665 1560 1845 1575
rect 300 1530 435 1560
rect 615 1545 690 1560
rect 750 1545 810 1560
rect 945 1545 1005 1560
rect 1080 1545 1155 1560
rect 1275 1545 1350 1560
rect 1410 1545 1485 1560
rect 1650 1545 1860 1560
rect 2025 1545 2235 1575
rect 2430 1560 2535 1590
rect 630 1530 705 1545
rect 735 1530 795 1545
rect 960 1530 1035 1545
rect 1065 1530 1140 1545
rect 1290 1530 1365 1545
rect 1395 1530 1470 1545
rect 1620 1530 1845 1545
rect 2025 1530 2220 1545
rect 285 1515 435 1530
rect 645 1515 780 1530
rect 975 1515 1125 1530
rect 1305 1515 1455 1530
rect 1605 1515 1830 1530
rect 2025 1515 2205 1530
rect 270 1485 435 1515
rect 660 1500 765 1515
rect 990 1500 1110 1515
rect 1320 1500 1440 1515
rect 1590 1500 1815 1515
rect 2025 1500 2190 1515
rect 675 1485 750 1500
rect 255 1455 300 1485
rect 240 1425 285 1455
rect 225 1395 270 1425
rect 210 1380 255 1395
rect 195 1365 255 1380
rect 195 1335 240 1365
rect 180 1320 240 1335
rect 180 1290 225 1320
rect 315 1290 435 1485
rect 690 1470 765 1485
rect 1005 1470 1095 1500
rect 1335 1485 1425 1500
rect 1575 1485 1800 1500
rect 1335 1470 1410 1485
rect 1560 1470 1785 1485
rect 2025 1470 2175 1500
rect 705 1455 780 1470
rect 990 1455 1110 1470
rect 1320 1455 1395 1470
rect 1545 1455 1770 1470
rect 2025 1455 2160 1470
rect 720 1440 795 1455
rect 975 1440 1125 1455
rect 1305 1440 1380 1455
rect 1530 1440 1755 1455
rect 735 1425 795 1440
rect 960 1425 1035 1440
rect 1065 1425 1125 1440
rect 1290 1425 1365 1440
rect 1515 1425 1740 1440
rect 2025 1425 2145 1455
rect 750 1410 810 1425
rect 945 1410 1020 1425
rect 1080 1410 1140 1425
rect 1275 1410 1350 1425
rect 1500 1410 1725 1425
rect 2025 1410 2130 1425
rect 765 1395 840 1410
rect 930 1395 1005 1410
rect 1095 1395 1155 1410
rect 1260 1395 1335 1410
rect 1470 1395 1695 1410
rect 1785 1395 1815 1410
rect 2025 1395 2115 1410
rect 780 1380 855 1395
rect 915 1380 990 1395
rect 1110 1380 1170 1395
rect 1245 1380 1320 1395
rect 1455 1380 1680 1395
rect 1770 1380 1830 1395
rect 795 1365 870 1380
rect 900 1365 975 1380
rect 1125 1365 1185 1380
rect 1230 1365 1305 1380
rect 1440 1365 1665 1380
rect 1755 1365 1845 1380
rect 2025 1365 2100 1395
rect 810 1350 960 1365
rect 1140 1350 1290 1365
rect 1410 1350 1650 1365
rect 1740 1350 1860 1365
rect 2025 1350 2085 1365
rect 825 1335 945 1350
rect 1155 1335 1275 1350
rect 1395 1335 1620 1350
rect 1725 1335 1785 1350
rect 1800 1335 1875 1350
rect 2025 1335 2070 1350
rect 840 1320 930 1335
rect 1170 1320 1260 1335
rect 1380 1320 1605 1335
rect 1710 1320 1770 1335
rect 1815 1320 1890 1335
rect 2025 1320 2055 1335
rect 855 1305 915 1320
rect 1185 1305 1245 1320
rect 1350 1305 1590 1320
rect 1695 1305 1755 1320
rect 1830 1305 1905 1320
rect 2025 1305 2040 1320
rect 870 1290 885 1305
rect 1200 1290 1215 1305
rect 1335 1290 1560 1305
rect 1680 1290 1740 1305
rect 1860 1290 1920 1305
rect 165 1230 225 1290
rect 330 1260 435 1290
rect 1305 1275 1545 1290
rect 1665 1275 1725 1290
rect 1875 1275 1935 1290
rect 2430 1275 2550 1560
rect 1290 1260 1515 1275
rect 1650 1260 1710 1275
rect 1890 1260 1950 1275
rect 165 1170 210 1230
rect 330 1200 450 1260
rect 1260 1245 1500 1260
rect 1620 1245 1695 1260
rect 1905 1245 1965 1260
rect 2430 1245 2535 1275
rect 1245 1230 1470 1245
rect 1605 1230 1680 1245
rect 1215 1215 1455 1230
rect 1605 1215 1665 1230
rect 1200 1200 1440 1215
rect 1590 1200 1680 1215
rect 1920 1200 1980 1245
rect 345 1185 450 1200
rect 1170 1185 1410 1200
rect 1575 1185 1695 1200
rect 1905 1185 1965 1200
rect 2415 1185 2535 1245
rect 165 1110 225 1170
rect 345 1140 465 1185
rect 1155 1170 1380 1185
rect 1560 1170 1620 1185
rect 1635 1170 1710 1185
rect 1890 1170 1950 1185
rect 2415 1170 2520 1185
rect 1125 1155 1365 1170
rect 1545 1155 1605 1170
rect 1650 1155 1725 1170
rect 1875 1155 1935 1170
rect 1095 1140 1335 1155
rect 1530 1140 1590 1155
rect 1665 1140 1740 1155
rect 1860 1140 1920 1155
rect 360 1125 465 1140
rect 1080 1125 1305 1140
rect 1515 1125 1575 1140
rect 1680 1125 1755 1140
rect 1830 1125 1905 1140
rect 2400 1125 2520 1170
rect 165 1095 240 1110
rect 180 1080 240 1095
rect 360 1080 480 1125
rect 1050 1110 1275 1125
rect 1500 1110 1560 1125
rect 1695 1110 1770 1125
rect 1815 1110 1890 1125
rect 1020 1095 1260 1110
rect 1485 1095 1545 1110
rect 1710 1095 1785 1110
rect 1800 1095 1875 1110
rect 990 1080 1230 1095
rect 1470 1080 1530 1095
rect 1725 1080 1860 1095
rect 2385 1080 2505 1125
rect 180 1065 255 1080
rect 180 1050 270 1065
rect 195 1035 270 1050
rect 375 1050 495 1080
rect 960 1065 1200 1080
rect 1455 1065 1515 1080
rect 1740 1065 1845 1080
rect 930 1050 1170 1065
rect 1440 1050 1500 1065
rect 1755 1050 1830 1065
rect 375 1035 510 1050
rect 900 1035 1140 1050
rect 1440 1035 1515 1050
rect 1740 1035 1845 1050
rect 2370 1035 2490 1080
rect 210 1020 300 1035
rect 420 1020 510 1035
rect 855 1020 1110 1035
rect 1455 1020 1530 1035
rect 1725 1020 1860 1035
rect 210 1005 315 1020
rect 480 1005 510 1020
rect 825 1005 1080 1020
rect 1470 1005 1545 1020
rect 1725 1005 1785 1020
rect 1800 1005 1875 1020
rect 2355 1005 2475 1035
rect 225 990 330 1005
rect 780 990 1050 1005
rect 1485 990 1560 1005
rect 1710 990 1770 1005
rect 1815 990 1890 1005
rect 2340 990 2475 1005
rect 240 975 360 990
rect 735 975 1020 990
rect 1500 975 1575 990
rect 1695 975 1755 990
rect 1830 975 1905 990
rect 2340 975 2460 990
rect 255 960 405 975
rect 690 960 975 975
rect 1515 960 1590 975
rect 1680 960 1740 975
rect 1845 960 1920 975
rect 2325 960 2460 975
rect 285 945 480 960
rect 600 945 945 960
rect 1530 945 1605 960
rect 1665 945 1725 960
rect 1860 945 1935 960
rect 2325 945 2445 960
rect 300 930 900 945
rect 1545 930 1620 945
rect 1650 930 1710 945
rect 1875 930 1950 945
rect 2310 930 2445 945
rect 330 915 855 930
rect 1560 915 1695 930
rect 1890 915 1965 930
rect 2310 915 2430 930
rect 360 900 810 915
rect 1575 900 1680 915
rect 1905 900 1980 915
rect 390 885 750 900
rect 1590 885 1665 900
rect 465 870 675 885
rect 1590 870 1680 885
rect 1920 870 1980 900
rect 2295 900 2430 915
rect 2295 885 2415 900
rect 2280 870 2415 885
rect 1575 855 1695 870
rect 1905 855 1965 870
rect 1560 840 1620 855
rect 1635 840 1710 855
rect 1890 840 1950 855
rect 2265 840 2400 870
rect 2640 855 2655 870
rect 2625 840 2655 855
rect 1545 825 1605 840
rect 1650 825 1725 840
rect 1875 825 1935 840
rect 2250 825 2385 840
rect 1530 810 1590 825
rect 1665 810 1740 825
rect 1860 810 1920 825
rect 2235 810 2370 825
rect 2625 810 2670 840
rect 495 795 645 810
rect 1515 795 1575 810
rect 1680 795 1755 810
rect 1845 795 1905 810
rect 2220 795 2370 810
rect 2610 795 2685 810
rect 510 780 660 795
rect 1500 780 1560 795
rect 1695 780 1770 795
rect 1830 780 1890 795
rect 2220 780 2355 795
rect 2595 780 2700 795
rect 525 765 660 780
rect 1485 765 1545 780
rect 1710 765 1785 780
rect 1815 765 1875 780
rect 2205 765 2340 780
rect 2580 765 2715 780
rect 525 750 675 765
rect 1470 750 1530 765
rect 1725 750 1860 765
rect 2190 750 2340 765
rect 2550 750 2745 765
rect 540 735 690 750
rect 1455 735 1515 750
rect 1740 735 1845 750
rect 2175 735 2325 750
rect 2520 735 2775 750
rect 555 720 705 735
rect 1440 720 1500 735
rect 1755 720 1830 735
rect 2160 720 2310 735
rect 2565 720 2730 735
rect 570 705 720 720
rect 1440 705 1515 720
rect 1755 705 1815 720
rect 2145 705 2295 720
rect 2580 705 2700 720
rect 585 690 735 705
rect 1455 690 1530 705
rect 1740 690 1800 705
rect 2130 690 2295 705
rect 2595 690 2685 705
rect 600 675 750 690
rect 1470 675 1545 690
rect 1725 675 1785 690
rect 2115 675 2280 690
rect 2610 675 2670 690
rect 600 660 765 675
rect 1485 660 1560 675
rect 1710 660 1770 675
rect 2100 660 2265 675
rect 2625 660 2670 675
rect 630 645 780 660
rect 1500 645 1575 660
rect 1695 645 1755 660
rect 2085 645 2250 660
rect 2625 645 2655 660
rect 645 630 810 645
rect 1515 630 1590 645
rect 1680 630 1740 645
rect 2070 630 2235 645
rect 2640 630 2655 645
rect 660 615 825 630
rect 1530 615 1605 630
rect 1665 615 1725 630
rect 2040 615 2220 630
rect 660 600 840 615
rect 1545 600 1605 615
rect 1650 600 1710 615
rect 2025 600 2205 615
rect 675 585 870 600
rect 1560 585 1695 600
rect 2010 585 2190 600
rect 705 570 885 585
rect 1575 570 1680 585
rect 1980 570 2175 585
rect 720 555 915 570
rect 1590 555 1665 570
rect 1965 555 2145 570
rect 735 540 930 555
rect 1605 540 1650 555
rect 1935 540 2130 555
rect 750 525 960 540
rect 1905 525 2115 540
rect 780 510 990 525
rect 1875 510 2100 525
rect 795 495 1020 510
rect 1845 495 2070 510
rect 810 480 1065 495
rect 1800 480 2055 495
rect 840 465 1095 480
rect 1770 465 2025 480
rect 870 450 1155 465
rect 1725 450 1995 465
rect 900 435 1200 450
rect 1665 435 1980 450
rect 915 420 1290 435
rect 1575 420 1950 435
rect 945 405 1920 420
rect 975 390 1890 405
rect 1005 375 1860 390
rect 1050 360 1815 375
rect 1095 345 1770 360
rect 1155 330 1710 345
rect 1215 315 1650 330
rect 1320 300 1545 315
<< fillblock >>
rect 0 0 2865 2865
<< properties >>
string FIXED_BBOX 0 0 2865 2865
string GDS_END 91846
string GDS_FILE ../../gds/gf180mcu_ws_ip__logo.gds
string GDS_START 114
<< end >>
