magic
tech gf180mcuD
magscale 1 10
timestamp 1766090161
<< metal1 >>
rect 464621 150317 465655 150325
rect 464621 150294 467095 150317
rect 464621 150087 464682 150294
rect 465587 150197 467095 150294
rect 465587 150087 465655 150197
rect 464621 150031 465655 150087
rect 464630 149669 465664 149707
rect 464630 149462 464699 149669
rect 465604 149533 465664 149669
rect 465604 149462 467095 149533
rect 464630 149413 467095 149462
rect 179939 87784 181643 88084
rect 179988 85019 180475 85319
rect 181343 85102 181643 87784
rect 180175 80199 180475 85019
rect 182534 84918 186777 85152
rect 187353 84918 187426 85152
rect 182050 80199 182350 80917
rect 180175 79899 182350 80199
<< via1 >>
rect 464682 150087 465587 150294
rect 324899 149906 325589 149997
rect 464699 149462 465604 149669
rect 324895 149125 325585 149216
rect 186777 84918 187353 85152
rect 128540 75303 128595 75355
rect 101868 75205 101923 75257
rect 102740 75205 102795 75257
rect 127668 75205 127723 75257
<< metal2 >>
rect 102880 292525 102956 430844
rect 128680 294553 128756 430844
rect 154480 296702 154556 430844
rect 180280 297381 180356 430844
rect 180280 297305 244161 297381
rect 154480 296626 243482 296702
rect 128680 294477 241333 294553
rect 102880 292449 239305 292525
rect 239229 232525 239305 292449
rect 241257 234553 241333 294477
rect 243406 236702 243482 296626
rect 244085 237381 244161 297305
rect 257680 239772 257756 430844
rect 283480 242154 283556 430844
rect 309280 243440 309356 430844
rect 309280 243364 322709 243440
rect 283480 242078 320709 242154
rect 257680 239696 318709 239772
rect 244085 237305 316709 237381
rect 243406 236626 314709 236702
rect 241257 234477 312709 234553
rect 239229 232449 310709 232525
rect 87550 136828 87650 175928
rect 87932 137028 88032 232328
rect 89052 146692 89128 204128
rect 310633 150752 310709 232449
rect 312633 150752 312709 234477
rect 314633 150752 314709 236626
rect 316633 150752 316709 237305
rect 318633 150752 318709 239696
rect 320633 150752 320709 242078
rect 322633 150752 322709 243364
rect 335080 209577 335156 430847
rect 360880 417502 360956 430793
rect 386680 419370 386756 430781
rect 412480 420911 412556 430789
rect 412480 420835 437030 420911
rect 386680 419294 435287 419370
rect 360880 417426 433959 417502
rect 324633 209501 335156 209577
rect 324633 150752 324709 209501
rect 433883 204920 433959 417426
rect 435211 205666 435287 419294
rect 436954 206527 437030 420835
rect 438280 207451 438356 430781
rect 464080 208407 464156 430789
rect 489880 420080 489956 430802
rect 468714 420004 489956 420080
rect 468714 209689 468790 420004
rect 515680 418225 515756 430796
rect 470575 418149 515756 418225
rect 470575 210624 470651 418149
rect 541480 416603 541556 430786
rect 619172 428709 619248 430801
rect 644972 429124 645048 430780
rect 670772 429613 670848 430785
rect 696572 430085 696648 430844
rect 471732 416527 541556 416603
rect 471732 211496 471808 416527
rect 471732 211420 482533 211496
rect 470575 210548 480533 210624
rect 468714 209613 478533 209689
rect 464080 208331 476533 208407
rect 438280 207375 474533 207451
rect 436954 206451 472533 206527
rect 435211 205590 470533 205666
rect 433883 204844 468533 204920
rect 468457 151343 468533 204844
rect 470457 151343 470533 205590
rect 472457 151343 472533 206451
rect 474457 151343 474533 207375
rect 476457 151343 476533 208331
rect 478457 151343 478533 209613
rect 480457 151343 480533 210548
rect 482457 151343 482533 211420
rect 463415 150294 465647 150328
rect 463415 150286 464682 150294
rect 89752 75169 89828 146528
rect 121870 142822 122027 147777
rect 122583 141216 122740 147777
rect 123332 138813 123488 147777
rect 128639 139024 128795 147777
rect 129110 143007 129267 147777
rect 129388 141423 129545 147777
rect 129703 141631 129860 147777
rect 129983 143214 130140 147777
rect 130454 139224 130611 147777
rect 136161 139427 136318 147777
rect 136948 141827 137105 147777
rect 137222 143419 137379 147777
rect 140121 146425 140278 147777
rect 140496 146632 140653 147790
rect 140870 146012 141027 147777
rect 141359 145812 141516 147777
rect 142167 144833 142324 147777
rect 143352 144633 143509 147777
rect 144536 144426 144692 147777
rect 148977 146239 149134 147777
rect 115552 75169 115628 75510
rect 154772 75426 154848 146328
rect 155805 141038 155962 147777
rect 158206 145624 158363 147777
rect 158657 145425 158814 147777
rect 159180 145239 159337 147777
rect 159951 145040 160108 147777
rect 163378 143630 163535 147777
rect 163846 142028 164003 147777
rect 164436 139622 164593 147777
rect 169942 139821 170099 147777
rect 170413 143843 170570 147777
rect 170692 142241 170848 147777
rect 171207 142441 171363 147777
rect 171487 144022 171643 147777
rect 171958 140021 172114 147777
rect 177664 140220 177821 147777
rect 178252 142633 178409 147777
rect 178726 144215 178883 147777
rect 246438 142815 246595 147848
rect 247151 141239 247308 147848
rect 247900 137224 248056 147848
rect 253207 137418 253363 147848
rect 253678 143019 253835 147848
rect 253956 141415 254113 147848
rect 254271 141614 254428 147848
rect 254551 143224 254708 147848
rect 255022 137631 255179 147848
rect 186777 87078 187353 87226
rect 180249 86247 180832 86303
rect 180776 80526 180832 86247
rect 186777 85192 187353 86550
rect 186743 85152 187391 85192
rect 186743 84918 186777 85152
rect 187353 84918 187391 85152
rect 186743 84887 187391 84918
rect 186777 84545 187353 84887
rect 181800 80526 181856 80710
rect 180776 80470 181856 80526
rect 182359 78593 182415 80994
rect 180291 78537 182415 78593
rect 180291 75384 180347 78537
rect 257972 75425 258048 145928
rect 260729 137816 260886 147848
rect 261516 141819 261673 147848
rect 261790 143430 261947 147848
rect 264689 146426 264846 147848
rect 265438 146021 265595 147848
rect 265927 145829 266084 147848
rect 266735 144815 266892 147848
rect 267920 144603 268077 147848
rect 269104 144424 269260 147848
rect 273545 146227 273702 147848
rect 280373 140830 280530 147848
rect 282774 145618 282931 147848
rect 283225 145426 283382 147848
rect 283748 145215 283905 147848
rect 284519 145023 284676 147848
rect 285869 131296 285945 145728
rect 287946 143622 288103 147848
rect 288414 142017 288571 147848
rect 289004 138019 289161 147848
rect 294510 138211 294667 147848
rect 294981 143827 295138 147848
rect 295260 142228 295416 147848
rect 295775 142446 295931 147848
rect 296055 144032 296211 147848
rect 296526 138416 296682 147848
rect 302232 138601 302389 147848
rect 302820 142598 302977 147848
rect 303294 144230 303451 147848
rect 308267 137028 308343 150241
rect 463415 150087 463488 150286
rect 464497 150087 464682 150286
rect 465587 150087 465647 150294
rect 463415 150031 465647 150087
rect 324882 150015 326730 150021
rect 324882 149997 325977 150015
rect 324882 149906 324899 149997
rect 325589 149921 325977 149997
rect 326701 149921 326730 150015
rect 325589 149906 326730 149921
rect 324882 149892 326730 149906
rect 463427 149669 465659 149711
rect 463427 149470 463492 149669
rect 464501 149470 464699 149669
rect 463427 149462 464699 149470
rect 465604 149462 465659 149669
rect 463427 149414 465659 149462
rect 324877 149216 326725 149234
rect 324877 149125 324895 149216
rect 325585 149210 326725 149216
rect 325585 149125 325964 149210
rect 324877 149116 325964 149125
rect 326688 149116 326725 149210
rect 324877 149105 326725 149116
rect 310217 148127 310282 148795
rect 310721 148277 310786 148795
rect 310721 148212 310953 148277
rect 310217 148062 310709 148127
rect 283772 131220 285945 131296
rect 283772 75356 283848 131220
rect 309572 75418 309648 145528
rect 310633 137202 310709 148062
rect 310888 148072 310953 148212
rect 311633 148072 311709 148073
rect 310888 148007 311709 148072
rect 311633 138814 311709 148007
rect 312121 148065 312186 148795
rect 312625 148218 312690 148795
rect 312625 148153 313016 148218
rect 312121 148000 312709 148065
rect 312633 137426 312709 148000
rect 312951 148058 313016 148153
rect 312951 147993 313709 148058
rect 313633 138992 313709 147993
rect 314025 148047 314090 148795
rect 314529 148277 314594 148795
rect 314529 148212 314971 148277
rect 314906 148065 314971 148212
rect 315929 148076 315994 148795
rect 316433 148255 316498 148795
rect 316433 148190 317273 148255
rect 317208 148083 317273 148190
rect 314025 147982 314709 148047
rect 314906 148000 315709 148065
rect 315929 148011 316709 148076
rect 317208 148018 317709 148083
rect 314633 137616 314709 147982
rect 315633 139197 315709 148000
rect 316633 137799 316709 148011
rect 317633 139395 317709 148018
rect 317833 148056 317898 148795
rect 318337 148242 318402 148795
rect 319737 148478 319802 148795
rect 319737 148413 319950 148478
rect 318337 148177 319709 148242
rect 317833 147991 318709 148056
rect 319632 148039 319709 148177
rect 318633 138034 318709 147991
rect 319633 139586 319709 148039
rect 319885 148085 319950 148413
rect 320241 148215 320306 148795
rect 321641 148275 321706 148795
rect 320241 148150 320989 148215
rect 321641 148210 321950 148275
rect 319885 148020 320709 148085
rect 320633 138217 320709 148020
rect 320924 148039 320989 148150
rect 321885 148041 321950 148210
rect 322145 148253 322210 148795
rect 323545 148271 323610 148795
rect 324049 148478 324114 148795
rect 324049 148413 324309 148478
rect 322145 148188 322999 148253
rect 323545 148206 323947 148271
rect 320924 147974 321709 148039
rect 321885 147976 322709 148041
rect 321633 139791 321709 147974
rect 322633 138413 322709 147976
rect 322934 148034 322999 148188
rect 323882 148058 323947 148206
rect 324244 148268 324309 148413
rect 324244 148203 325709 148268
rect 322934 147969 323709 148034
rect 323882 147993 324709 148058
rect 323633 140022 323709 147969
rect 324633 138609 324709 147993
rect 325633 140220 325709 148203
rect 335372 75356 335448 145328
rect 361172 75356 361248 145128
rect 386972 75355 387048 144928
rect 412772 75356 412848 144728
rect 438572 75352 438648 144504
rect 464372 75356 464448 144328
rect 465840 136840 465916 150561
rect 468041 147985 468106 149084
rect 468545 148135 468610 149084
rect 468545 148070 468777 148135
rect 468041 147920 468533 147985
rect 468457 137203 468533 147920
rect 468712 147930 468777 148070
rect 469457 147930 469533 147931
rect 468712 147865 469533 147930
rect 469457 138804 469533 147865
rect 469945 147923 470010 149084
rect 470449 148076 470514 149084
rect 470449 148011 470840 148076
rect 469945 147858 470533 147923
rect 470457 137432 470533 147858
rect 470775 147916 470840 148011
rect 470775 147851 471533 147916
rect 471457 139007 471533 147851
rect 471849 147905 471914 149084
rect 472353 148135 472418 149084
rect 472353 148070 472795 148135
rect 472730 147923 472795 148070
rect 473753 147934 473818 149084
rect 474257 148113 474322 149084
rect 474257 148048 475097 148113
rect 475032 147941 475097 148048
rect 471849 147840 472533 147905
rect 472730 147858 473533 147923
rect 473753 147869 474533 147934
rect 475032 147876 475533 147941
rect 472457 137615 472533 147840
rect 473457 139210 473533 147858
rect 474457 137824 474533 147869
rect 475457 139433 475533 147876
rect 475657 147914 475722 149084
rect 476161 148100 476226 149084
rect 477561 148336 477626 149084
rect 477561 148271 477774 148336
rect 476161 148035 477533 148100
rect 475657 147849 476533 147914
rect 477456 147897 477533 148035
rect 476457 138014 476533 147849
rect 477457 139629 477533 147897
rect 477709 147943 477774 148271
rect 478065 148073 478130 149084
rect 479465 148133 479530 149084
rect 478065 148008 478813 148073
rect 479465 148068 479774 148133
rect 477709 147878 478533 147943
rect 478457 138216 478533 147878
rect 478748 147897 478813 148008
rect 479709 147899 479774 148068
rect 479969 148111 480034 149084
rect 481369 148129 481434 149084
rect 481873 148336 481938 149084
rect 481873 148271 482133 148336
rect 479969 148046 480823 148111
rect 481369 148064 481771 148129
rect 478748 147832 479533 147897
rect 479709 147834 480533 147899
rect 479457 139838 479533 147832
rect 480457 138406 480533 147834
rect 480758 147892 480823 148046
rect 481706 147916 481771 148064
rect 482068 148126 482133 148271
rect 482068 148061 483533 148126
rect 480758 147827 481533 147892
rect 481706 147851 482533 147916
rect 481457 140014 481533 147827
rect 482457 138629 482533 147851
rect 483457 140230 483533 148061
rect 487071 142832 487228 147281
rect 487784 141251 487941 147281
rect 488533 138838 488689 147281
rect 490172 75356 490248 144128
rect 493840 139017 493996 147281
rect 494311 143033 494468 147281
rect 494589 141416 494746 147281
rect 494904 141625 495061 147281
rect 495184 143215 495341 147281
rect 495655 139206 495812 147281
rect 501362 139423 501519 147281
rect 502149 141829 502306 147281
rect 502423 143428 502580 147281
rect 505322 146425 505479 147281
rect 506559 145827 506717 147281
rect 507368 144826 507525 147281
rect 508553 144618 508710 147281
rect 509737 144430 509893 147281
rect 514178 146237 514335 147281
rect 515972 75356 516048 143928
rect 521006 140639 521163 147281
rect 523407 145612 523564 147281
rect 523858 145431 524015 147281
rect 524381 145223 524538 147281
rect 525152 145028 525309 147281
rect 528579 143616 528736 147281
rect 529047 142010 529204 147281
rect 529637 139625 529794 147281
rect 535143 139808 535300 147281
rect 535614 143809 535771 147281
rect 535893 142227 536049 147281
rect 536408 142428 536564 147281
rect 536688 144016 536844 147281
rect 537159 140009 537315 147281
rect 541772 75355 541848 143729
rect 542865 140197 543022 147281
rect 543453 142602 543610 147281
rect 543927 144204 544084 147281
rect 602627 142815 602784 147281
rect 603340 141212 603497 147281
rect 604089 137204 604245 147281
rect 609396 137421 609552 147281
rect 609867 143033 610024 147281
rect 610145 141429 610302 147281
rect 610460 141617 610617 147281
rect 610740 143221 610897 147281
rect 611211 137619 611368 147281
rect 616918 137809 617075 147281
rect 617705 141803 617862 147281
rect 617979 143414 618136 147281
rect 620878 146390 621035 147281
rect 622115 145809 622273 147281
rect 622924 144811 623081 147281
rect 624109 144589 624266 147281
rect 625293 144412 625449 147281
rect 629734 146219 629891 147281
rect 619172 75356 619248 143528
rect 636562 140433 636719 147281
rect 638963 145616 639120 147281
rect 639414 145408 639571 147281
rect 639937 145220 640094 147281
rect 640708 145022 640865 147281
rect 644135 143627 644292 147281
rect 644603 142003 644760 147281
rect 645193 138015 645350 147281
rect 646741 131258 646817 143328
rect 650699 138213 650856 147281
rect 651170 143805 651327 147281
rect 651449 142211 651605 147281
rect 651964 142409 652120 147281
rect 652244 144012 652400 147281
rect 652715 138421 652871 147281
rect 658421 138639 658578 147281
rect 659009 142617 659166 147281
rect 659483 144210 659640 147281
rect 644972 131182 646817 131258
rect 644972 75356 645048 131182
rect 670772 75356 670848 143128
rect 696572 75356 696648 142928
rect 697213 141031 697289 161156
rect 697907 140833 697983 189348
rect 698515 140644 698591 217543
rect 699167 140434 699243 245753
rect 699596 142642 699672 428786
rect 699996 142448 700072 429198
rect 700311 142239 700387 429692
rect 700668 142048 700744 430156
rect 701025 141843 701101 358551
rect 701404 141656 701480 330339
rect 701789 141433 701865 302147
rect 702157 141238 702233 273948
<< via2 >>
rect 186777 86550 187353 87078
rect 463488 150087 464497 150286
rect 325977 149921 326701 150015
rect 463492 149470 464501 149669
rect 325964 149116 326688 149210
<< metal3 >>
rect 696572 430077 700744 430153
rect 670682 429614 700387 429690
rect 644888 429124 700072 429199
rect 645100 429123 700072 429124
rect 619156 428710 699672 428786
rect 701027 358472 710913 358548
rect 701402 330272 710929 330348
rect 701763 302072 710912 302148
rect 702149 273872 710911 273948
rect 180778 249660 218272 250360
rect 220172 249660 220752 250360
rect 222802 249660 223122 250360
rect 225172 249660 225828 250360
rect 227878 249660 228198 250360
rect 230248 249660 230828 250360
rect 232655 249660 232910 250360
rect 180810 249071 192472 249581
rect 194372 249071 194952 249581
rect 197002 249071 197322 249581
rect 199372 249071 200028 249581
rect 202078 249071 202398 249581
rect 204448 249071 205028 249581
rect 206851 249071 232930 249581
rect 180810 248481 218272 248971
rect 220172 248481 220752 248971
rect 222802 248481 223122 248971
rect 225172 248481 225828 248971
rect 227878 248481 228198 248971
rect 230248 248481 230828 248971
rect 232655 248481 232930 248971
rect 180810 247859 192472 248369
rect 194372 247859 194952 248369
rect 197002 247859 197322 248369
rect 199372 247859 200028 248369
rect 202078 247859 202398 248369
rect 204448 247859 205028 248369
rect 206851 247859 232930 248369
rect 180810 247269 218272 247759
rect 220172 247269 220752 247759
rect 222802 247269 223122 247759
rect 225172 247269 225828 247759
rect 227878 247269 228198 247759
rect 230248 247269 230828 247759
rect 232655 247269 232930 247759
rect 180810 246647 192472 247157
rect 194372 246647 194952 247157
rect 197002 246647 197322 247157
rect 199372 246647 200028 247157
rect 202078 246647 202398 247157
rect 204448 246647 205028 247157
rect 206851 246647 232930 247157
rect 180810 246057 218272 246547
rect 220172 246057 220752 246547
rect 222802 246057 223122 246547
rect 225172 246057 225828 246547
rect 227878 246057 228198 246547
rect 230248 246057 230828 246547
rect 232655 246057 232930 246547
rect 180810 245435 192472 245945
rect 194372 245435 194952 245945
rect 197002 245435 197322 245945
rect 199372 245435 200028 245945
rect 202078 245435 202398 245945
rect 204448 245435 205028 245945
rect 206851 245435 232930 245945
rect 699087 245672 710900 245748
rect 180810 244845 218272 245335
rect 220172 244845 220752 245335
rect 222802 244845 223122 245335
rect 225172 244845 225828 245335
rect 227878 244845 228198 245335
rect 230248 244845 230828 245335
rect 232655 244845 232930 245335
rect 180810 244223 192472 244733
rect 194372 244223 194952 244733
rect 197002 244223 197322 244733
rect 199372 244223 200028 244733
rect 202078 244223 202398 244733
rect 204448 244223 205028 244733
rect 206851 244223 232930 244733
rect 180810 243633 218272 244123
rect 220172 243633 220752 244123
rect 222802 243633 223122 244123
rect 225172 243633 225828 244123
rect 227878 243633 228198 244123
rect 230248 243633 230828 244123
rect 232655 243633 232930 244123
rect 180810 243011 192472 243521
rect 194372 243011 194952 243521
rect 197002 243011 197322 243521
rect 199372 243011 200028 243521
rect 202078 243011 202398 243521
rect 204448 243011 205028 243521
rect 206851 243011 232930 243521
rect 180810 242421 218272 242911
rect 220172 242421 220752 242911
rect 222802 242421 223122 242911
rect 225172 242421 225828 242911
rect 227878 242421 228198 242911
rect 230248 242421 230828 242911
rect 232655 242421 232930 242911
rect 180810 241799 192472 242309
rect 194372 241799 194952 242309
rect 197002 241799 197322 242309
rect 199372 241799 200028 242309
rect 202078 241799 202398 242309
rect 204448 241799 205028 242309
rect 206851 241799 232930 242309
rect 180810 241209 218272 241699
rect 220172 241209 220752 241699
rect 222802 241209 223122 241699
rect 225172 241209 225828 241699
rect 227878 241209 228198 241699
rect 230248 241209 230828 241699
rect 232655 241209 232930 241699
rect 180810 240587 192472 241097
rect 194372 240587 194952 241097
rect 197002 240587 197322 241097
rect 199372 240587 200028 241097
rect 202078 240587 202398 241097
rect 204448 240587 205028 241097
rect 206851 240587 232930 241097
rect 180810 239997 218272 240487
rect 220172 239997 220752 240487
rect 222802 239997 223122 240487
rect 225172 239997 225828 240487
rect 227878 239997 228198 240487
rect 230248 239997 230828 240487
rect 232655 239997 232930 240487
rect 180810 239375 192472 239885
rect 194372 239375 194952 239885
rect 197002 239375 197322 239885
rect 199372 239375 200028 239885
rect 202078 239375 202398 239885
rect 204448 239375 205028 239885
rect 206851 239375 232930 239885
rect 180810 238785 218272 239275
rect 220172 238785 220752 239275
rect 222802 238785 223122 239275
rect 225172 238785 225828 239275
rect 227878 238785 228198 239275
rect 230248 238785 230828 239275
rect 232655 238785 232930 239275
rect 180810 238163 192472 238673
rect 194372 238163 194952 238673
rect 197002 238163 197322 238673
rect 199372 238163 200028 238673
rect 202078 238163 202398 238673
rect 204448 238163 205028 238673
rect 206851 238163 232930 238673
rect 180810 237573 218272 238063
rect 220172 237573 220752 238063
rect 222802 237573 223122 238063
rect 225172 237573 225828 238063
rect 227878 237573 228198 238063
rect 230248 237573 230828 238063
rect 232655 237573 232930 238063
rect 180810 236951 192472 237461
rect 194372 236951 194952 237461
rect 197002 236951 197322 237461
rect 199372 236951 200028 237461
rect 202078 236951 202398 237461
rect 204448 236951 205028 237461
rect 206851 236951 232930 237461
rect 180810 236361 218272 236851
rect 220172 236361 220752 236851
rect 222802 236361 223122 236851
rect 225172 236361 225828 236851
rect 227878 236361 228198 236851
rect 230248 236361 230828 236851
rect 232655 236361 232930 236851
rect 180810 235739 192472 236249
rect 194372 235739 194952 236249
rect 197002 235739 197322 236249
rect 199372 235739 200028 236249
rect 202078 235739 202398 236249
rect 204448 235739 205028 236249
rect 206851 235739 232930 236249
rect 180810 235149 218272 235639
rect 220172 235149 220752 235639
rect 222802 235149 223122 235639
rect 225172 235149 225828 235639
rect 227878 235149 228198 235639
rect 230248 235149 230828 235639
rect 232655 235149 232930 235639
rect 180810 234527 192472 235037
rect 194372 234527 194952 235037
rect 197002 234527 197322 235037
rect 199372 234527 200028 235037
rect 202078 234527 202398 235037
rect 204448 234527 205028 235037
rect 206851 234527 232930 235037
rect 180810 233937 218272 234427
rect 220172 233937 220752 234427
rect 222802 233937 223122 234427
rect 225172 233937 225828 234427
rect 227878 233937 228198 234427
rect 230248 233937 230828 234427
rect 232655 233937 232930 234427
rect 180810 233315 192472 233825
rect 194372 233315 194952 233825
rect 197002 233315 197322 233825
rect 199372 233315 200028 233825
rect 202078 233315 202398 233825
rect 204448 233315 205028 233825
rect 206851 233315 232930 233825
rect 180810 232725 218272 233215
rect 220172 232725 220752 233215
rect 222802 232725 223122 233215
rect 225172 232725 225828 233215
rect 227878 232725 228198 233215
rect 230248 232725 230828 233215
rect 232655 232725 232930 233215
rect 75470 232252 87932 232328
rect 180810 232103 192472 232613
rect 194372 232103 194952 232613
rect 197002 232103 197322 232613
rect 199372 232103 200028 232613
rect 202078 232103 202398 232613
rect 204448 232103 205028 232613
rect 206851 232103 232930 232613
rect 180810 231513 218272 232003
rect 220172 231513 220752 232003
rect 222802 231513 223122 232003
rect 225172 231513 225828 232003
rect 227878 231513 228198 232003
rect 230248 231513 230828 232003
rect 232655 231513 232930 232003
rect 180810 230891 192472 231401
rect 194372 230891 194952 231401
rect 197002 230891 197322 231401
rect 199372 230891 200028 231401
rect 202078 230891 202398 231401
rect 204448 230891 205028 231401
rect 206851 230891 232930 231401
rect 180810 230301 218272 230791
rect 220172 230301 220752 230791
rect 222802 230301 223122 230791
rect 225172 230301 225828 230791
rect 227878 230301 228198 230791
rect 230248 230301 230828 230791
rect 232655 230301 232930 230791
rect 180810 229679 192472 230189
rect 194372 229679 194952 230189
rect 197002 229679 197322 230189
rect 199372 229679 200028 230189
rect 202078 229679 202398 230189
rect 204448 229679 205028 230189
rect 206851 229679 232930 230189
rect 180810 229089 218272 229579
rect 220172 229089 220752 229579
rect 222802 229089 223122 229579
rect 225172 229089 225828 229579
rect 227878 229089 228198 229579
rect 230248 229089 230828 229579
rect 232655 229089 232930 229579
rect 180810 228467 192472 228977
rect 194372 228467 194952 228977
rect 197002 228467 197322 228977
rect 199372 228467 200028 228977
rect 202078 228467 202398 228977
rect 204448 228467 205028 228977
rect 206851 228467 232930 228977
rect 180810 227877 218272 228367
rect 220172 227877 220752 228367
rect 222802 227877 223122 228367
rect 225172 227877 225828 228367
rect 227878 227877 228198 228367
rect 230248 227877 230828 228367
rect 232655 227877 232930 228367
rect 180810 227255 192472 227765
rect 194372 227255 194952 227765
rect 197002 227255 197322 227765
rect 199372 227255 200028 227765
rect 202078 227255 202398 227765
rect 204448 227255 205028 227765
rect 206851 227255 232930 227765
rect 180810 226665 218272 227155
rect 220172 226665 220752 227155
rect 222802 226665 223122 227155
rect 225172 226665 225828 227155
rect 227878 226665 228198 227155
rect 230248 226665 230828 227155
rect 232655 226665 232930 227155
rect 180810 226043 192472 226553
rect 194372 226043 194952 226553
rect 197002 226043 197322 226553
rect 199372 226043 200028 226553
rect 202078 226043 202398 226553
rect 204448 226043 205028 226553
rect 206851 226043 232930 226553
rect 180810 225453 218272 225943
rect 220172 225453 220752 225943
rect 222802 225453 223122 225943
rect 225172 225453 225828 225943
rect 227878 225453 228198 225943
rect 230248 225453 230828 225943
rect 232655 225453 232930 225943
rect 180810 224831 192472 225341
rect 194372 224831 194952 225341
rect 197002 224831 197322 225341
rect 199372 224831 200028 225341
rect 202078 224831 202398 225341
rect 204448 224831 205028 225341
rect 206851 224831 232930 225341
rect 180810 224241 218272 224731
rect 220172 224241 220752 224731
rect 222802 224241 223122 224731
rect 225172 224241 225828 224731
rect 227878 224241 228198 224731
rect 230248 224241 230828 224731
rect 232655 224241 232930 224731
rect 180810 223619 192472 224129
rect 194372 223619 194952 224129
rect 197002 223619 197322 224129
rect 199372 223619 200028 224129
rect 202078 223619 202398 224129
rect 204448 223619 205028 224129
rect 206851 223619 232930 224129
rect 180810 223029 218272 223519
rect 220172 223029 220752 223519
rect 222802 223029 223122 223519
rect 225172 223029 225828 223519
rect 227878 223029 228198 223519
rect 230248 223029 230828 223519
rect 232655 223029 232930 223519
rect 180810 222407 192472 222917
rect 194372 222407 194952 222917
rect 197002 222407 197322 222917
rect 199372 222407 200028 222917
rect 202078 222407 202398 222917
rect 204448 222407 205028 222917
rect 206851 222407 232930 222917
rect 180810 221817 218272 222307
rect 220172 221817 220752 222307
rect 222802 221817 223122 222307
rect 225172 221817 225828 222307
rect 227878 221817 228198 222307
rect 230248 221817 230828 222307
rect 232655 221817 232930 222307
rect 180810 221195 192472 221705
rect 194372 221195 194952 221705
rect 197002 221195 197322 221705
rect 199372 221195 200028 221705
rect 202078 221195 202398 221705
rect 204448 221195 205028 221705
rect 206851 221195 232930 221705
rect 180810 220605 218272 221095
rect 220172 220605 220752 221095
rect 222802 220605 223122 221095
rect 225172 220605 225828 221095
rect 227878 220605 228198 221095
rect 230248 220605 230828 221095
rect 232655 220605 232930 221095
rect 180810 219983 192472 220493
rect 194372 219983 194952 220493
rect 197002 219983 197322 220493
rect 199372 219983 200028 220493
rect 202078 219983 202398 220493
rect 204448 219983 205028 220493
rect 206851 219983 232930 220493
rect 180810 219393 218272 219883
rect 220172 219393 220752 219883
rect 222802 219393 223122 219883
rect 225172 219393 225828 219883
rect 227878 219393 228198 219883
rect 230248 219393 230828 219883
rect 232655 219393 232930 219883
rect 180810 218771 192472 219281
rect 194372 218771 194952 219281
rect 197002 218771 197322 219281
rect 199372 218771 200028 219281
rect 202078 218771 202398 219281
rect 204448 218771 205028 219281
rect 206851 218771 232930 219281
rect 180810 218181 218272 218671
rect 220172 218181 220752 218671
rect 222802 218181 223122 218671
rect 225172 218181 225828 218671
rect 227878 218181 228198 218671
rect 230248 218181 230828 218671
rect 232655 218181 232930 218671
rect 180810 217559 192472 218069
rect 194372 217559 194952 218069
rect 197002 217559 197322 218069
rect 199372 217559 200028 218069
rect 202078 217559 202398 218069
rect 204448 217559 205028 218069
rect 206851 217559 232930 218069
rect 698436 217472 710903 217548
rect 180810 216969 218272 217459
rect 220172 216969 220752 217459
rect 222802 216969 223122 217459
rect 225172 216969 225828 217459
rect 227878 216969 228198 217459
rect 230248 216969 230828 217459
rect 232655 216969 232930 217459
rect 180810 216347 192472 216857
rect 194372 216347 194952 216857
rect 197002 216347 197322 216857
rect 199372 216347 200028 216857
rect 202078 216347 202398 216857
rect 204448 216347 205028 216857
rect 206851 216347 232930 216857
rect 180810 215757 218272 216247
rect 220172 215757 220752 216247
rect 222802 215757 223122 216247
rect 225172 215757 225828 216247
rect 227878 215757 228198 216247
rect 230248 215757 230828 216247
rect 232655 215757 232930 216247
rect 180810 215135 192472 215645
rect 194372 215135 194952 215645
rect 197002 215135 197322 215645
rect 199372 215135 200028 215645
rect 202078 215135 202398 215645
rect 204448 215135 205028 215645
rect 206851 215135 232930 215645
rect 180810 214545 218272 215035
rect 220172 214545 220752 215035
rect 222802 214545 223122 215035
rect 225172 214545 225828 215035
rect 227878 214545 228198 215035
rect 230248 214545 230828 215035
rect 232655 214545 232930 215035
rect 180810 213923 192472 214433
rect 194372 213923 194952 214433
rect 197002 213923 197322 214433
rect 199372 213923 200028 214433
rect 202078 213923 202398 214433
rect 204448 213923 205028 214433
rect 206851 213923 232930 214433
rect 180810 213333 218272 213823
rect 220172 213333 220752 213823
rect 222802 213333 223122 213823
rect 225172 213333 225828 213823
rect 227878 213333 228198 213823
rect 230248 213333 230828 213823
rect 232655 213333 232930 213823
rect 180810 212711 192472 213221
rect 194372 212711 194952 213221
rect 197002 212711 197322 213221
rect 199372 212711 200028 213221
rect 202078 212711 202398 213221
rect 204448 212711 205028 213221
rect 206851 212711 232930 213221
rect 180810 212121 218272 212611
rect 220172 212121 220752 212611
rect 222802 212121 223122 212611
rect 225172 212121 225828 212611
rect 227878 212121 228198 212611
rect 230248 212121 230828 212611
rect 232655 212121 232930 212611
rect 180810 211499 192472 212009
rect 194372 211499 194952 212009
rect 197002 211499 197322 212009
rect 199372 211499 200028 212009
rect 202078 211499 202398 212009
rect 204448 211499 205028 212009
rect 206851 211499 206950 212009
rect 218180 211399 218272 211576
rect 180810 210909 218272 211399
rect 218180 210876 218272 210909
rect 220172 210876 220752 211576
rect 222802 210876 223122 211576
rect 225172 210876 225828 211576
rect 227878 210876 228198 211576
rect 230248 210876 230828 211576
rect 232655 210876 245202 211576
rect 180778 210287 192472 210797
rect 194372 210287 194952 210797
rect 197002 210287 197322 210797
rect 199372 210287 200028 210797
rect 202078 210287 202398 210797
rect 204448 210287 205028 210797
rect 206851 210287 245202 210797
rect 180778 209697 218272 210187
rect 220172 209697 220752 210187
rect 222802 209697 223122 210187
rect 225172 209697 225828 210187
rect 227878 209697 228198 210187
rect 230248 209697 230828 210187
rect 232655 209697 245202 210187
rect 180778 209095 192472 209585
rect 194372 209095 194952 209585
rect 197002 209095 197322 209585
rect 199372 209095 200028 209585
rect 202078 209095 202398 209585
rect 204448 209095 205028 209585
rect 206851 209095 245202 209585
rect 180778 208485 218272 208975
rect 220172 208485 220752 208975
rect 222802 208485 223122 208975
rect 225172 208485 225828 208975
rect 227878 208485 228198 208975
rect 230248 208485 230828 208975
rect 232655 208485 245202 208975
rect 180778 207883 192472 208373
rect 194372 207883 194952 208373
rect 197002 207883 197322 208373
rect 199372 207883 200028 208373
rect 202078 207883 202398 208373
rect 204448 207883 205028 208373
rect 206851 207883 245202 208373
rect 180778 207273 218272 207763
rect 220172 207273 220752 207763
rect 222802 207273 223122 207763
rect 225172 207273 225828 207763
rect 227878 207273 228198 207763
rect 230248 207273 230828 207763
rect 232655 207273 245202 207763
rect 180778 206671 192472 207161
rect 194372 206671 194952 207161
rect 197002 206671 197322 207161
rect 199372 206671 200028 207161
rect 202078 206671 202398 207161
rect 204448 206671 205028 207161
rect 206851 206671 245202 207161
rect 180778 206061 218272 206551
rect 220172 206061 220752 206551
rect 222802 206061 223122 206551
rect 225172 206061 225828 206551
rect 227878 206061 228198 206551
rect 230248 206061 230828 206551
rect 232655 206061 245202 206551
rect 180778 205459 192472 205949
rect 194372 205459 194952 205949
rect 197002 205459 197322 205949
rect 199372 205459 200028 205949
rect 202078 205459 202398 205949
rect 204448 205459 205028 205949
rect 206851 205459 245202 205949
rect 180778 204849 218272 205339
rect 220172 204849 220752 205339
rect 222802 204849 223122 205339
rect 225172 204849 225828 205339
rect 227878 204849 228198 205339
rect 230248 204849 230828 205339
rect 232655 204849 245202 205339
rect 180778 204247 192472 204737
rect 194372 204247 194952 204737
rect 197002 204247 197322 204737
rect 199372 204247 200028 204737
rect 202078 204247 202398 204737
rect 204448 204247 205028 204737
rect 206851 204247 245202 204737
rect 75390 204052 89128 204128
rect 180778 203637 218272 204127
rect 220172 203637 220752 204127
rect 222802 203637 223122 204127
rect 225172 203637 225828 204127
rect 227878 203637 228198 204127
rect 230248 203637 230828 204127
rect 232655 203637 245202 204127
rect 180778 203035 192472 203525
rect 194372 203035 194952 203525
rect 197002 203035 197322 203525
rect 199372 203035 200028 203525
rect 202078 203035 202398 203525
rect 204448 203035 205028 203525
rect 206851 203035 245202 203525
rect 180778 202425 218272 202915
rect 220172 202425 220752 202915
rect 222802 202425 223122 202915
rect 225172 202425 225828 202915
rect 227878 202425 228198 202915
rect 230248 202425 230828 202915
rect 232655 202425 245202 202915
rect 180778 201823 192472 202313
rect 194372 201823 194952 202313
rect 197002 201823 197322 202313
rect 199372 201823 200028 202313
rect 202078 201823 202398 202313
rect 204448 201823 205028 202313
rect 206851 201823 245202 202313
rect 180778 201213 218272 201703
rect 220172 201213 220752 201703
rect 222802 201213 223122 201703
rect 225172 201213 225828 201703
rect 227878 201213 228198 201703
rect 230248 201213 230828 201703
rect 232655 201213 245202 201703
rect 180778 200611 192472 201101
rect 194372 200611 194952 201101
rect 197002 200611 197322 201101
rect 199372 200611 200028 201101
rect 202078 200611 202398 201101
rect 204448 200611 205028 201101
rect 206851 200611 245202 201101
rect 180778 200001 218272 200491
rect 220172 200001 220752 200491
rect 222802 200001 223122 200491
rect 225172 200001 225828 200491
rect 227878 200001 228198 200491
rect 230248 200001 230828 200491
rect 232655 200001 245202 200491
rect 180778 199399 192472 199889
rect 194372 199399 194952 199889
rect 197002 199399 197322 199889
rect 199372 199399 200028 199889
rect 202078 199399 202398 199889
rect 204448 199399 205028 199889
rect 206851 199399 245202 199889
rect 180778 198789 218272 199279
rect 220172 198789 220752 199279
rect 222802 198789 223122 199279
rect 225172 198789 225828 199279
rect 227878 198789 228198 199279
rect 230248 198789 230828 199279
rect 232655 198789 245202 199279
rect 180778 198187 192472 198677
rect 194372 198187 194952 198677
rect 197002 198187 197322 198677
rect 199372 198187 200028 198677
rect 202078 198187 202398 198677
rect 204448 198187 205028 198677
rect 206851 198187 245202 198677
rect 180778 197577 218272 198067
rect 220172 197577 220752 198067
rect 222802 197577 223122 198067
rect 225172 197577 225828 198067
rect 227878 197577 228198 198067
rect 230248 197577 230828 198067
rect 232655 197577 245202 198067
rect 180778 196975 192472 197465
rect 194372 196975 194952 197465
rect 197002 196975 197322 197465
rect 199372 196975 200028 197465
rect 202078 196975 202398 197465
rect 204448 196975 205028 197465
rect 206851 196975 245202 197465
rect 180778 196365 218272 196855
rect 220172 196365 220752 196855
rect 222802 196365 223122 196855
rect 225172 196365 225828 196855
rect 227878 196365 228198 196855
rect 230248 196365 230828 196855
rect 232655 196365 245202 196855
rect 180778 195763 192472 196253
rect 194372 195763 194952 196253
rect 197002 195763 197322 196253
rect 199372 195763 200028 196253
rect 202078 195763 202398 196253
rect 204448 195763 205028 196253
rect 206851 195763 245202 196253
rect 180778 195153 218272 195643
rect 220172 195153 220752 195643
rect 222802 195153 223122 195643
rect 225172 195153 225828 195643
rect 227878 195153 228198 195643
rect 230248 195153 230828 195643
rect 232655 195153 245202 195643
rect 180778 194551 192472 195041
rect 194372 194551 194952 195041
rect 197002 194551 197322 195041
rect 199372 194551 200028 195041
rect 202078 194551 202398 195041
rect 204448 194551 205028 195041
rect 206851 194551 245202 195041
rect 180778 193941 218272 194431
rect 220172 193941 220752 194431
rect 222802 193941 223122 194431
rect 225172 193941 225828 194431
rect 227878 193941 228198 194431
rect 230248 193941 230828 194431
rect 232655 193941 245202 194431
rect 180778 193339 192472 193829
rect 194372 193339 194952 193829
rect 197002 193339 197322 193829
rect 199372 193339 200028 193829
rect 202078 193339 202398 193829
rect 204448 193339 205028 193829
rect 206851 193339 245202 193829
rect 180778 192729 218272 193219
rect 220172 192729 220752 193219
rect 222802 192729 223122 193219
rect 225172 192729 225828 193219
rect 227878 192729 228198 193219
rect 230248 192729 230828 193219
rect 232655 192729 245202 193219
rect 180778 192127 192472 192617
rect 194372 192127 194952 192617
rect 197002 192127 197322 192617
rect 199372 192127 200028 192617
rect 202078 192127 202398 192617
rect 204448 192127 205028 192617
rect 206851 192127 245202 192617
rect 180778 191517 218272 192007
rect 220172 191517 220752 192007
rect 222802 191517 223122 192007
rect 225172 191517 225828 192007
rect 227878 191517 228198 192007
rect 230248 191517 230828 192007
rect 232655 191517 245202 192007
rect 180778 190915 192472 191405
rect 194372 190915 194952 191405
rect 197002 190915 197322 191405
rect 199372 190915 200028 191405
rect 202078 190915 202398 191405
rect 204448 190915 205028 191405
rect 206851 190915 245202 191405
rect 545982 190983 579472 191683
rect 581372 190983 581952 191683
rect 584002 190983 584322 191683
rect 586372 190983 587028 191683
rect 589078 190983 589398 191683
rect 591448 190983 592028 191683
rect 593928 190983 601325 191683
rect 180778 190305 218272 190795
rect 220172 190305 220752 190795
rect 222802 190305 223122 190795
rect 225172 190305 225828 190795
rect 227878 190305 228198 190795
rect 230248 190305 230828 190795
rect 232655 190305 245202 190795
rect 545982 190394 553672 190904
rect 555572 190394 556152 190904
rect 558202 190394 558522 190904
rect 560572 190394 561228 190904
rect 563278 190394 563598 190904
rect 565648 190394 566228 190904
rect 568128 190394 601325 190904
rect 180778 189703 192472 190193
rect 194372 189703 194952 190193
rect 197002 189703 197322 190193
rect 199372 189703 200028 190193
rect 202078 189703 202398 190193
rect 204448 189703 205028 190193
rect 206851 189703 245202 190193
rect 545982 189804 579472 190294
rect 581372 189804 581952 190294
rect 584002 189804 584322 190294
rect 586372 189804 587028 190294
rect 589078 189804 589398 190294
rect 591448 189804 592028 190294
rect 593928 189804 601325 190294
rect 180778 189093 218272 189583
rect 220172 189093 220752 189583
rect 222802 189093 223122 189583
rect 225172 189093 225828 189583
rect 227878 189093 228198 189583
rect 230248 189093 230828 189583
rect 232655 189093 245202 189583
rect 545982 189202 553672 189692
rect 555572 189202 556152 189692
rect 558202 189202 558522 189692
rect 560572 189202 561228 189692
rect 563278 189202 563598 189692
rect 565648 189202 566228 189692
rect 568128 189202 601325 189692
rect 697842 189272 710912 189348
rect 180778 188491 192472 188981
rect 194372 188491 194952 188981
rect 197002 188491 197322 188981
rect 199372 188491 200028 188981
rect 202078 188491 202398 188981
rect 204448 188491 205028 188981
rect 206851 188491 245202 188981
rect 545982 188592 579472 189082
rect 581372 188592 581952 189082
rect 584002 188592 584322 189082
rect 586372 188592 587028 189082
rect 589078 188592 589398 189082
rect 591448 188592 592028 189082
rect 593928 188592 601325 189082
rect 180778 187881 218272 188371
rect 220172 187881 220752 188371
rect 222802 187881 223122 188371
rect 225172 187881 225828 188371
rect 227878 187881 228198 188371
rect 230248 187881 230828 188371
rect 232655 187881 245202 188371
rect 545982 187990 553672 188480
rect 555572 187990 556152 188480
rect 558202 187990 558522 188480
rect 560572 187990 561228 188480
rect 563278 187990 563598 188480
rect 565648 187990 566228 188480
rect 568128 187990 601325 188480
rect 180778 187279 192472 187769
rect 194372 187279 194952 187769
rect 197002 187279 197322 187769
rect 199372 187279 200028 187769
rect 202078 187279 202398 187769
rect 204448 187279 205028 187769
rect 206851 187279 245202 187769
rect 545982 187380 579472 187870
rect 581372 187380 581952 187870
rect 584002 187380 584322 187870
rect 586372 187380 587028 187870
rect 589078 187380 589398 187870
rect 591448 187380 592028 187870
rect 593928 187380 601325 187870
rect 180778 186669 218272 187159
rect 220172 186669 220752 187159
rect 222802 186669 223122 187159
rect 225172 186669 225828 187159
rect 227878 186669 228198 187159
rect 230248 186669 230828 187159
rect 232655 186669 245202 187159
rect 545982 186778 553672 187268
rect 555572 186778 556152 187268
rect 558202 186778 558522 187268
rect 560572 186778 561228 187268
rect 563278 186778 563598 187268
rect 565648 186778 566228 187268
rect 568128 186778 601325 187268
rect 180778 186067 192472 186557
rect 194372 186067 194952 186557
rect 197002 186067 197322 186557
rect 199372 186067 200028 186557
rect 202078 186067 202398 186557
rect 204448 186067 205028 186557
rect 206851 186067 245202 186557
rect 545982 186168 579472 186658
rect 581372 186168 581952 186658
rect 584002 186168 584322 186658
rect 586372 186168 587028 186658
rect 589078 186168 589398 186658
rect 591448 186168 592028 186658
rect 593928 186168 601325 186658
rect 180778 185457 218272 185947
rect 220172 185457 220752 185947
rect 222802 185457 223122 185947
rect 225172 185457 225828 185947
rect 227878 185457 228198 185947
rect 230248 185457 230828 185947
rect 232655 185457 245202 185947
rect 545982 185566 553672 186056
rect 555572 185566 556152 186056
rect 558202 185566 558522 186056
rect 560572 185566 561228 186056
rect 563278 185566 563598 186056
rect 565648 185566 566228 186056
rect 568128 185566 601325 186056
rect 180778 184855 192472 185345
rect 194372 184855 194952 185345
rect 197002 184855 197322 185345
rect 199372 184855 200028 185345
rect 202078 184855 202398 185345
rect 204448 184855 205028 185345
rect 206851 184855 245202 185345
rect 545982 184956 579472 185446
rect 581372 184956 581952 185446
rect 584002 184956 584322 185446
rect 586372 184956 587028 185446
rect 589078 184956 589398 185446
rect 591448 184956 592028 185446
rect 593928 184956 601325 185446
rect 180778 184245 218272 184735
rect 220172 184245 220752 184735
rect 222802 184245 223122 184735
rect 225172 184245 225828 184735
rect 227878 184245 228198 184735
rect 230248 184245 230828 184735
rect 232655 184245 245202 184735
rect 545982 184354 553672 184844
rect 555572 184354 556152 184844
rect 558202 184354 558522 184844
rect 560572 184354 561228 184844
rect 563278 184354 563598 184844
rect 565648 184354 566228 184844
rect 568128 184354 601325 184844
rect 180778 183643 192472 184133
rect 194372 183643 194952 184133
rect 197002 183643 197322 184133
rect 199372 183643 200028 184133
rect 202078 183643 202398 184133
rect 204448 183643 205028 184133
rect 206851 183643 245202 184133
rect 545982 183744 579472 184234
rect 581372 183744 581952 184234
rect 584002 183744 584322 184234
rect 586372 183744 587028 184234
rect 589078 183744 589398 184234
rect 591448 183744 592028 184234
rect 593928 183744 601325 184234
rect 180778 183033 218272 183523
rect 220172 183033 220752 183523
rect 222802 183033 223122 183523
rect 225172 183033 225828 183523
rect 227878 183033 228198 183523
rect 230248 183033 230828 183523
rect 232655 183033 245202 183523
rect 545982 183142 553672 183632
rect 555572 183142 556152 183632
rect 558202 183142 558522 183632
rect 560572 183142 561228 183632
rect 563278 183142 563598 183632
rect 565648 183142 566228 183632
rect 568128 183142 601325 183632
rect 180778 182431 192472 182921
rect 194372 182431 194952 182921
rect 197002 182431 197322 182921
rect 199372 182431 200028 182921
rect 202078 182431 202398 182921
rect 204448 182431 205028 182921
rect 206851 182431 245202 182921
rect 545982 182532 579472 183022
rect 581372 182532 581952 183022
rect 584002 182532 584322 183022
rect 586372 182532 587028 183022
rect 589078 182532 589398 183022
rect 591448 182532 592028 183022
rect 593928 182532 601325 183022
rect 180778 181821 218272 182311
rect 220172 181821 220752 182311
rect 222802 181821 223122 182311
rect 225172 181821 225828 182311
rect 227878 181821 228198 182311
rect 230248 181821 230828 182311
rect 232655 181821 245202 182311
rect 545982 181930 553672 182420
rect 555572 181930 556152 182420
rect 558202 181930 558522 182420
rect 560572 181930 561228 182420
rect 563278 181930 563598 182420
rect 565648 181930 566228 182420
rect 568128 181930 601325 182420
rect 180778 181219 192472 181709
rect 194372 181219 194952 181709
rect 197002 181219 197322 181709
rect 199372 181219 200028 181709
rect 202078 181219 202398 181709
rect 204448 181219 205028 181709
rect 206851 181219 245202 181709
rect 545982 181320 579472 181810
rect 581372 181320 581952 181810
rect 584002 181320 584322 181810
rect 586372 181320 587028 181810
rect 589078 181320 589398 181810
rect 591448 181320 592028 181810
rect 593928 181320 601325 181810
rect 180778 180609 218272 181099
rect 220172 180609 220752 181099
rect 222802 180609 223122 181099
rect 225172 180609 225828 181099
rect 227878 180609 228198 181099
rect 230248 180609 230828 181099
rect 232655 180609 245202 181099
rect 545982 180718 553672 181208
rect 555572 180718 556152 181208
rect 558202 180718 558522 181208
rect 560572 180718 561228 181208
rect 563278 180718 563598 181208
rect 565648 180718 566228 181208
rect 568128 180718 601325 181208
rect 180778 180007 192472 180497
rect 194372 180007 194952 180497
rect 197002 180007 197322 180497
rect 199372 180007 200028 180497
rect 202078 180007 202398 180497
rect 204448 180007 205028 180497
rect 206851 180007 245202 180497
rect 545982 180108 579472 180598
rect 581372 180108 581952 180598
rect 584002 180108 584322 180598
rect 586372 180108 587028 180598
rect 589078 180108 589398 180598
rect 591448 180108 592028 180598
rect 593928 180108 601325 180598
rect 180778 179397 218272 179887
rect 220172 179397 220752 179887
rect 222802 179397 223122 179887
rect 225172 179397 225828 179887
rect 227878 179397 228198 179887
rect 230248 179397 230828 179887
rect 232655 179397 245202 179887
rect 545982 179506 553672 179996
rect 555572 179506 556152 179996
rect 558202 179506 558522 179996
rect 560572 179506 561228 179996
rect 563278 179506 563598 179996
rect 565648 179506 566228 179996
rect 568128 179506 601325 179996
rect 180778 178795 192472 179285
rect 194372 178795 194952 179285
rect 197002 178795 197322 179285
rect 199372 178795 200028 179285
rect 202078 178795 202398 179285
rect 204448 178795 205028 179285
rect 206851 178795 245202 179285
rect 545982 178896 579472 179386
rect 581372 178896 581952 179386
rect 584002 178896 584322 179386
rect 586372 178896 587028 179386
rect 589078 178896 589398 179386
rect 591448 178896 592028 179386
rect 593928 178896 601325 179386
rect 180778 178185 218272 178675
rect 220172 178185 220752 178675
rect 222802 178185 223122 178675
rect 225172 178185 225828 178675
rect 227878 178185 228198 178675
rect 230248 178185 230828 178675
rect 232655 178185 245202 178675
rect 545982 178294 553672 178784
rect 555572 178294 556152 178784
rect 558202 178294 558522 178784
rect 560572 178294 561228 178784
rect 563278 178294 563598 178784
rect 565648 178294 566228 178784
rect 568128 178294 601325 178784
rect 180778 177583 192472 178073
rect 194372 177583 194952 178073
rect 197002 177583 197322 178073
rect 199372 177583 200028 178073
rect 202078 177583 202398 178073
rect 204448 177583 205028 178073
rect 206851 177583 245202 178073
rect 545982 177684 579472 178174
rect 581372 177684 581952 178174
rect 584002 177684 584322 178174
rect 586372 177684 587028 178174
rect 589078 177684 589398 178174
rect 591448 177684 592028 178174
rect 593928 177684 601325 178174
rect 180778 176973 218272 177463
rect 220172 176973 220752 177463
rect 222802 176973 223122 177463
rect 225172 176973 225828 177463
rect 227878 176973 228198 177463
rect 230248 176973 230828 177463
rect 232655 176973 245202 177463
rect 545982 177082 553672 177572
rect 555572 177082 556152 177572
rect 558202 177082 558522 177572
rect 560572 177082 561228 177572
rect 563278 177082 563598 177572
rect 565648 177082 566228 177572
rect 568128 177082 601325 177572
rect 180778 176371 192472 176861
rect 194372 176371 194952 176861
rect 197002 176371 197322 176861
rect 199372 176371 200028 176861
rect 202078 176371 202398 176861
rect 204448 176371 205028 176861
rect 206851 176371 245202 176861
rect 545982 176472 579472 176962
rect 581372 176472 581952 176962
rect 584002 176472 584322 176962
rect 586372 176472 587028 176962
rect 589078 176472 589398 176962
rect 591448 176472 592028 176962
rect 593928 176472 601325 176962
rect 75465 175852 87550 175928
rect 180778 175761 218272 176251
rect 220172 175761 220752 176251
rect 222802 175761 223122 176251
rect 225172 175761 225828 176251
rect 227878 175761 228198 176251
rect 230248 175761 230828 176251
rect 232655 175761 245202 176251
rect 545982 175870 553672 176360
rect 555572 175870 556152 176360
rect 558202 175870 558522 176360
rect 560572 175870 561228 176360
rect 563278 175870 563598 176360
rect 565648 175870 566228 176360
rect 568128 175870 601325 176360
rect 180778 175159 192472 175649
rect 194372 175159 194952 175649
rect 197002 175159 197322 175649
rect 199372 175159 200028 175649
rect 202078 175159 202398 175649
rect 204448 175159 205028 175649
rect 206851 175159 245202 175649
rect 545982 175260 579472 175750
rect 581372 175260 581952 175750
rect 584002 175260 584322 175750
rect 586372 175260 587028 175750
rect 589078 175260 589398 175750
rect 591448 175260 592028 175750
rect 593928 175260 601325 175750
rect 180778 174549 218272 175039
rect 220172 174549 220752 175039
rect 222802 174549 223122 175039
rect 225172 174549 225828 175039
rect 227878 174549 228198 175039
rect 230248 174549 230828 175039
rect 232655 174549 245202 175039
rect 545982 174658 553672 175148
rect 555572 174658 556152 175148
rect 558202 174658 558522 175148
rect 560572 174658 561228 175148
rect 563278 174658 563598 175148
rect 565648 174658 566228 175148
rect 568128 174658 601325 175148
rect 180778 173947 192472 174437
rect 194372 173947 194952 174437
rect 197002 173947 197322 174437
rect 199372 173947 200028 174437
rect 202078 173947 202398 174437
rect 204448 173947 205028 174437
rect 206851 173947 245202 174437
rect 545982 174048 579472 174538
rect 581372 174048 581952 174538
rect 584002 174048 584322 174538
rect 586372 174048 587028 174538
rect 589078 174048 589398 174538
rect 591448 174048 592028 174538
rect 593928 174048 601325 174538
rect 180778 173337 218272 173827
rect 220172 173337 220752 173827
rect 222802 173337 223122 173827
rect 225172 173337 225828 173827
rect 227878 173337 228198 173827
rect 230248 173337 230828 173827
rect 232655 173337 245202 173827
rect 545982 173446 553672 173936
rect 555572 173446 556152 173936
rect 558202 173446 558522 173936
rect 560572 173446 561228 173936
rect 563278 173446 563598 173936
rect 565648 173446 566228 173936
rect 568128 173446 601325 173936
rect 180778 172735 192472 173225
rect 194372 172735 194952 173225
rect 197002 172735 197322 173225
rect 199372 172735 200028 173225
rect 202078 172735 202398 173225
rect 204448 172735 205028 173225
rect 206851 172735 245202 173225
rect 545982 172836 579472 173326
rect 581372 172836 581952 173326
rect 584002 172836 584322 173326
rect 586372 172836 587028 173326
rect 589078 172836 589398 173326
rect 591448 172836 592028 173326
rect 593928 172836 601325 173326
rect 180778 172125 218272 172615
rect 220172 172125 220752 172615
rect 222802 172125 223122 172615
rect 225172 172125 225828 172615
rect 227878 172125 228198 172615
rect 230248 172125 230828 172615
rect 232655 172125 245202 172615
rect 545982 172234 553672 172724
rect 555572 172234 556152 172724
rect 558202 172234 558522 172724
rect 560572 172234 561228 172724
rect 563278 172234 563598 172724
rect 565648 172234 566228 172724
rect 568128 172234 601325 172724
rect 180778 171523 192472 172013
rect 194372 171523 194952 172013
rect 197002 171523 197322 172013
rect 199372 171523 200028 172013
rect 202078 171523 202398 172013
rect 204448 171523 205028 172013
rect 206851 171523 245202 172013
rect 545982 171624 579472 172114
rect 581372 171624 581952 172114
rect 584002 171624 584322 172114
rect 586372 171624 587028 172114
rect 589078 171624 589398 172114
rect 591448 171624 592028 172114
rect 593928 171624 601325 172114
rect 180778 170913 218272 171403
rect 220172 170913 220752 171403
rect 222802 170913 223122 171403
rect 225172 170913 225828 171403
rect 227878 170913 228198 171403
rect 230248 170913 230828 171403
rect 232655 170913 245202 171403
rect 545982 171022 553672 171512
rect 555572 171022 556152 171512
rect 558202 171022 558522 171512
rect 560572 171022 561228 171512
rect 563278 171022 563598 171512
rect 565648 171022 566228 171512
rect 568128 171022 601325 171512
rect 180778 170027 192472 170630
rect 194372 170027 194952 170630
rect 197002 170027 197322 170630
rect 199372 170027 200028 170630
rect 202078 170027 202398 170630
rect 204448 170027 205028 170630
rect 206851 170027 245202 170630
rect 545982 170412 579472 170902
rect 581372 170412 581952 170902
rect 584002 170412 584322 170902
rect 586372 170412 587028 170902
rect 589078 170412 589398 170902
rect 591448 170412 592028 170902
rect 593928 170412 601325 170902
rect 180778 166792 218272 169740
rect 220172 166792 220752 169740
rect 222802 166792 223122 169740
rect 225172 166792 225828 169740
rect 227878 166792 228198 169740
rect 230248 166792 230828 169740
rect 232655 166792 245202 169740
rect 545982 169526 553672 170129
rect 555572 169526 556152 170129
rect 558202 169526 558522 170129
rect 560572 169526 561228 170129
rect 563278 169526 563598 170129
rect 565648 169526 566228 170129
rect 568128 169526 601325 170129
rect 180778 165136 192472 166524
rect 194372 165136 194952 166524
rect 197002 165136 197322 166524
rect 199372 165136 200028 166524
rect 202078 165136 202398 166524
rect 204448 165136 205028 166524
rect 206851 165136 245202 166524
rect 545982 166291 579472 169239
rect 581372 166291 581952 169239
rect 584002 166291 584322 169239
rect 586372 166291 587028 169239
rect 589078 166291 589398 169239
rect 591448 166291 592028 169239
rect 593928 166291 601325 169239
rect 545982 164635 553672 166023
rect 555572 164635 556152 166023
rect 558202 164635 558522 166023
rect 560572 164635 561228 166023
rect 563278 164635 563598 166023
rect 565648 164635 566228 166023
rect 568128 164635 601325 166023
rect 180778 162728 218272 163429
rect 220172 162728 220752 163429
rect 222802 162728 223122 163429
rect 225172 162728 225828 163429
rect 227878 162728 228198 163429
rect 230248 162728 230828 163429
rect 232655 162728 245202 163429
rect 180778 161629 192472 162330
rect 194372 161629 194952 162330
rect 197002 161629 197322 162330
rect 199372 161629 200028 162330
rect 202078 161629 202398 162330
rect 204448 161629 205028 162330
rect 206851 161629 245202 162330
rect 545982 162227 579472 162928
rect 581372 162227 581952 162928
rect 584002 162227 584322 162928
rect 586372 162227 587028 162928
rect 589078 162227 589398 162928
rect 591448 162227 592028 162928
rect 593928 162227 601325 162928
rect 180778 159399 218272 161308
rect 220172 159399 220752 161308
rect 222802 159399 223122 161308
rect 225172 159399 225828 161308
rect 227878 159399 228198 161308
rect 230248 159399 230828 161308
rect 232655 159399 245202 161308
rect 545982 161128 553672 161829
rect 555572 161128 556152 161829
rect 558202 161128 558522 161829
rect 560572 161128 561228 161829
rect 563278 161128 563598 161829
rect 565648 161128 566228 161829
rect 568128 161128 601325 161829
rect 697136 161072 710906 161148
rect 180778 157348 192472 159200
rect 194372 157348 194952 159200
rect 197002 157348 197322 159200
rect 199372 157348 200028 159200
rect 202078 157348 202398 159200
rect 204448 157348 205028 159200
rect 206851 157348 245202 159200
rect 545982 158898 579472 160807
rect 581372 158898 581952 160807
rect 584002 158898 584322 160807
rect 586372 158898 587028 160807
rect 589078 158898 589398 160807
rect 591448 158898 592028 160807
rect 593928 158898 601325 160807
rect 180778 155760 218272 157222
rect 220172 155760 220752 157222
rect 222802 155760 223122 157222
rect 225172 155760 225828 157222
rect 227878 155760 228198 157222
rect 230248 155760 230828 157222
rect 232655 155760 245202 157222
rect 545982 156847 553672 158699
rect 555572 156847 556152 158699
rect 558202 156847 558522 158699
rect 560572 156847 561228 158699
rect 563278 156847 563598 158699
rect 565648 156847 566228 158699
rect 568128 156847 601325 158699
rect 180778 154481 192472 155404
rect 194372 154481 194952 155404
rect 197002 154481 197322 155404
rect 199372 154481 200028 155404
rect 202078 154481 202398 155404
rect 204448 154481 205028 155404
rect 206851 154481 245202 155404
rect 545982 155259 579472 156721
rect 581372 155259 581952 156721
rect 584002 155259 584322 156721
rect 586372 155259 587028 156721
rect 589078 155259 589398 156721
rect 591448 155259 592028 156721
rect 593928 155259 601325 156721
rect 180778 153063 218272 154018
rect 220172 153063 220752 154018
rect 222802 153063 223122 154018
rect 225172 153063 225828 154018
rect 227878 153063 228198 154018
rect 230248 153063 230828 154018
rect 232655 153063 245202 154018
rect 545982 153980 553672 154903
rect 555572 153980 556152 154903
rect 558202 153980 558522 154903
rect 560572 153980 561228 154903
rect 563278 153980 563598 154903
rect 565648 153980 566228 154903
rect 568128 153980 601325 154903
rect 180778 151720 192472 152851
rect 194372 151720 194952 152851
rect 197002 151720 197322 152851
rect 199372 151720 200028 152851
rect 202078 151720 202398 152851
rect 204448 151720 205028 152851
rect 206851 151720 245202 152851
rect 545982 152562 579472 153517
rect 581372 152562 581952 153517
rect 584002 152562 584322 153517
rect 586372 152562 587028 153517
rect 589078 152562 589398 153517
rect 591448 152562 592028 153517
rect 593928 152562 601325 153517
rect 180778 150599 218272 151628
rect 220172 150599 220752 151628
rect 222802 150599 223122 151628
rect 225172 150599 225828 151628
rect 227878 150599 228198 151628
rect 230248 150599 230828 151628
rect 232655 150599 245202 151628
rect 545982 151219 553672 152350
rect 555572 151219 556152 152350
rect 558202 151219 558522 152350
rect 560572 151219 561228 152350
rect 563278 151219 563598 152350
rect 565648 151219 566228 152350
rect 568128 151219 601325 152350
rect 465826 150464 467068 150540
rect 180778 149508 192472 150397
rect 194372 149508 194952 150397
rect 197002 149508 197322 150397
rect 199372 149508 200028 150397
rect 202078 149508 202398 150397
rect 204448 149508 205028 150397
rect 206851 149508 245202 150397
rect 308151 150160 309264 150236
rect 459340 150035 459446 150332
rect 460246 150286 464573 150332
rect 460246 150087 463488 150286
rect 464497 150087 464573 150286
rect 545982 150098 579472 151127
rect 581372 150098 581952 151127
rect 584002 150098 584322 151127
rect 586372 150098 587028 151127
rect 589078 150098 589398 151127
rect 591448 150098 592028 151127
rect 593928 150098 601325 151127
rect 460246 150035 464573 150087
rect 325956 150015 328649 150030
rect 325956 149921 325977 150015
rect 326701 149921 328649 150015
rect 325956 149896 328649 149921
rect 329463 149896 329483 150030
rect 459366 149414 460979 149711
rect 461779 149669 464560 149711
rect 461779 149470 463492 149669
rect 464501 149470 464560 149669
rect 461779 149414 464560 149470
rect 180778 148620 218272 149320
rect 220172 148620 220752 149320
rect 222802 148620 223122 149320
rect 225172 148620 225828 149320
rect 227878 148620 228198 149320
rect 230248 148620 230828 149320
rect 232655 148620 245202 149320
rect 325931 149210 327021 149232
rect 325931 149116 325964 149210
rect 326688 149116 327021 149210
rect 325931 149098 327021 149116
rect 327835 149098 329458 149232
rect 545982 149007 553672 149896
rect 555572 149007 556152 149896
rect 558202 149007 558522 149896
rect 560572 149007 561228 149896
rect 563278 149007 563598 149896
rect 565648 149007 566228 149896
rect 568128 149007 601325 149896
rect 545982 148119 579472 148819
rect 581372 148119 581952 148819
rect 584002 148119 584322 148819
rect 586372 148119 587028 148819
rect 589078 148119 589398 148819
rect 591448 148119 592028 148819
rect 593928 148119 601325 148819
rect 75251 147639 78033 147739
rect 77933 146128 78033 147639
rect 89030 146628 140690 146728
rect 89752 146428 621112 146528
rect 120404 146228 630049 146328
rect 77933 146028 325936 146128
rect 120404 145828 622323 145928
rect 120404 145628 639215 145728
rect 120404 145428 639682 145528
rect 120404 145228 640202 145328
rect 120404 145028 640975 145128
rect 120404 144828 623158 144928
rect 120404 144628 624336 144728
rect 120404 144428 625550 144528
rect 120404 144228 659737 144328
rect 120404 144028 652551 144128
rect 120404 143828 651392 143928
rect 120404 143628 644402 143728
rect 120404 143428 619384 143528
rect 120404 143228 646945 143328
rect 120404 143028 671001 143128
rect 120404 142828 696808 142928
rect 120404 142628 699810 142728
rect 120404 142428 700187 142528
rect 120404 142228 700514 142328
rect 120404 142028 700586 142128
rect 120404 141828 701227 141928
rect 120404 141628 701612 141728
rect 120404 141428 701998 141528
rect 120404 141228 702365 141328
rect 155004 141028 697455 141128
rect 279604 140828 697998 140928
rect 520204 140628 698577 140728
rect 635804 140428 699344 140528
rect 120404 140228 325888 140328
rect 466986 140228 543137 140328
rect 120404 140028 323888 140128
rect 466986 140028 537421 140128
rect 120404 139828 321889 139928
rect 466986 139828 535386 139928
rect 120404 139628 319876 139728
rect 466988 139628 529882 139728
rect 120404 139428 317889 139528
rect 466986 139428 501588 139528
rect 120404 139228 315817 139328
rect 466986 139228 495895 139328
rect 120404 139028 313817 139128
rect 466986 139028 494077 139128
rect 120404 138828 311844 138928
rect 466986 138828 488809 138928
rect 245604 138628 324811 138728
rect 466986 138628 658722 138728
rect 245604 138428 322836 138528
rect 466996 138428 653011 138528
rect 245604 138228 320856 138328
rect 466990 138228 650953 138328
rect 245604 138028 318849 138128
rect 466990 138028 645440 138128
rect 245604 137828 316857 137928
rect 466986 137828 617175 137928
rect 245604 137628 314847 137728
rect 466986 137628 611500 137728
rect 245604 137428 312863 137528
rect 466986 137428 609694 137528
rect 245604 137228 310839 137328
rect 466981 137228 604350 137328
rect 88032 137028 308485 137128
rect 87650 136828 466072 136928
rect 186496 86550 186777 87078
rect 187353 86550 218272 87078
rect 220172 86550 220293 87078
<< via3 >>
rect 218272 249660 220172 250360
rect 220752 249660 222802 250360
rect 223122 249660 225172 250360
rect 225828 249660 227878 250360
rect 228198 249660 230248 250360
rect 230828 249660 232655 250360
rect 192472 249071 194372 249581
rect 194952 249071 197002 249581
rect 197322 249071 199372 249581
rect 200028 249071 202078 249581
rect 202398 249071 204448 249581
rect 205028 249071 206851 249581
rect 218272 248481 220172 248971
rect 220752 248481 222802 248971
rect 223122 248481 225172 248971
rect 225828 248481 227878 248971
rect 228198 248481 230248 248971
rect 230828 248481 232655 248971
rect 192472 247859 194372 248369
rect 194952 247859 197002 248369
rect 197322 247859 199372 248369
rect 200028 247859 202078 248369
rect 202398 247859 204448 248369
rect 205028 247859 206851 248369
rect 218272 247269 220172 247759
rect 220752 247269 222802 247759
rect 223122 247269 225172 247759
rect 225828 247269 227878 247759
rect 228198 247269 230248 247759
rect 230828 247269 232655 247759
rect 192472 246647 194372 247157
rect 194952 246647 197002 247157
rect 197322 246647 199372 247157
rect 200028 246647 202078 247157
rect 202398 246647 204448 247157
rect 205028 246647 206851 247157
rect 218272 246057 220172 246547
rect 220752 246057 222802 246547
rect 223122 246057 225172 246547
rect 225828 246057 227878 246547
rect 228198 246057 230248 246547
rect 230828 246057 232655 246547
rect 192472 245435 194372 245945
rect 194952 245435 197002 245945
rect 197322 245435 199372 245945
rect 200028 245435 202078 245945
rect 202398 245435 204448 245945
rect 205028 245435 206851 245945
rect 75272 245239 75332 245298
rect 218272 244845 220172 245335
rect 220752 244845 222802 245335
rect 223122 244845 225172 245335
rect 225828 244845 227878 245335
rect 228198 244845 230248 245335
rect 230828 244845 232655 245335
rect 75272 244367 75332 244426
rect 192472 244223 194372 244733
rect 194952 244223 197002 244733
rect 197322 244223 199372 244733
rect 200028 244223 202078 244733
rect 202398 244223 204448 244733
rect 205028 244223 206851 244733
rect 218272 243633 220172 244123
rect 220752 243633 222802 244123
rect 223122 243633 225172 244123
rect 225828 243633 227878 244123
rect 228198 243633 230248 244123
rect 230828 243633 232655 244123
rect 192472 243011 194372 243521
rect 194952 243011 197002 243521
rect 197322 243011 199372 243521
rect 200028 243011 202078 243521
rect 202398 243011 204448 243521
rect 205028 243011 206851 243521
rect 218272 242421 220172 242911
rect 220752 242421 222802 242911
rect 223122 242421 225172 242911
rect 225828 242421 227878 242911
rect 228198 242421 230248 242911
rect 230828 242421 232655 242911
rect 192472 241799 194372 242309
rect 194952 241799 197002 242309
rect 197322 241799 199372 242309
rect 200028 241799 202078 242309
rect 202398 241799 204448 242309
rect 205028 241799 206851 242309
rect 218272 241209 220172 241699
rect 220752 241209 222802 241699
rect 223122 241209 225172 241699
rect 225828 241209 227878 241699
rect 228198 241209 230248 241699
rect 230828 241209 232655 241699
rect 192472 240587 194372 241097
rect 194952 240587 197002 241097
rect 197322 240587 199372 241097
rect 200028 240587 202078 241097
rect 202398 240587 204448 241097
rect 205028 240587 206851 241097
rect 218272 239997 220172 240487
rect 220752 239997 222802 240487
rect 223122 239997 225172 240487
rect 225828 239997 227878 240487
rect 228198 239997 230248 240487
rect 230828 239997 232655 240487
rect 192472 239375 194372 239885
rect 194952 239375 197002 239885
rect 197322 239375 199372 239885
rect 200028 239375 202078 239885
rect 202398 239375 204448 239885
rect 205028 239375 206851 239885
rect 218272 238785 220172 239275
rect 220752 238785 222802 239275
rect 223122 238785 225172 239275
rect 225828 238785 227878 239275
rect 228198 238785 230248 239275
rect 230828 238785 232655 239275
rect 192472 238163 194372 238673
rect 194952 238163 197002 238673
rect 197322 238163 199372 238673
rect 200028 238163 202078 238673
rect 202398 238163 204448 238673
rect 205028 238163 206851 238673
rect 218272 237573 220172 238063
rect 220752 237573 222802 238063
rect 223122 237573 225172 238063
rect 225828 237573 227878 238063
rect 228198 237573 230248 238063
rect 230828 237573 232655 238063
rect 192472 236951 194372 237461
rect 194952 236951 197002 237461
rect 197322 236951 199372 237461
rect 200028 236951 202078 237461
rect 202398 236951 204448 237461
rect 205028 236951 206851 237461
rect 218272 236361 220172 236851
rect 220752 236361 222802 236851
rect 223122 236361 225172 236851
rect 225828 236361 227878 236851
rect 228198 236361 230248 236851
rect 230828 236361 232655 236851
rect 192472 235739 194372 236249
rect 194952 235739 197002 236249
rect 197322 235739 199372 236249
rect 200028 235739 202078 236249
rect 202398 235739 204448 236249
rect 205028 235739 206851 236249
rect 218272 235149 220172 235639
rect 220752 235149 222802 235639
rect 223122 235149 225172 235639
rect 225828 235149 227878 235639
rect 228198 235149 230248 235639
rect 230828 235149 232655 235639
rect 192472 234527 194372 235037
rect 194952 234527 197002 235037
rect 197322 234527 199372 235037
rect 200028 234527 202078 235037
rect 202398 234527 204448 235037
rect 205028 234527 206851 235037
rect 218272 233937 220172 234427
rect 220752 233937 222802 234427
rect 223122 233937 225172 234427
rect 225828 233937 227878 234427
rect 228198 233937 230248 234427
rect 230828 233937 232655 234427
rect 192472 233315 194372 233825
rect 194952 233315 197002 233825
rect 197322 233315 199372 233825
rect 200028 233315 202078 233825
rect 202398 233315 204448 233825
rect 205028 233315 206851 233825
rect 218272 232725 220172 233215
rect 220752 232725 222802 233215
rect 223122 232725 225172 233215
rect 225828 232725 227878 233215
rect 228198 232725 230248 233215
rect 230828 232725 232655 233215
rect 192472 232103 194372 232613
rect 194952 232103 197002 232613
rect 197322 232103 199372 232613
rect 200028 232103 202078 232613
rect 202398 232103 204448 232613
rect 205028 232103 206851 232613
rect 218272 231513 220172 232003
rect 220752 231513 222802 232003
rect 223122 231513 225172 232003
rect 225828 231513 227878 232003
rect 228198 231513 230248 232003
rect 230828 231513 232655 232003
rect 192472 230891 194372 231401
rect 194952 230891 197002 231401
rect 197322 230891 199372 231401
rect 200028 230891 202078 231401
rect 202398 230891 204448 231401
rect 205028 230891 206851 231401
rect 218272 230301 220172 230791
rect 220752 230301 222802 230791
rect 223122 230301 225172 230791
rect 225828 230301 227878 230791
rect 228198 230301 230248 230791
rect 230828 230301 232655 230791
rect 192472 229679 194372 230189
rect 194952 229679 197002 230189
rect 197322 229679 199372 230189
rect 200028 229679 202078 230189
rect 202398 229679 204448 230189
rect 205028 229679 206851 230189
rect 218272 229089 220172 229579
rect 220752 229089 222802 229579
rect 223122 229089 225172 229579
rect 225828 229089 227878 229579
rect 228198 229089 230248 229579
rect 230828 229089 232655 229579
rect 192472 228467 194372 228977
rect 194952 228467 197002 228977
rect 197322 228467 199372 228977
rect 200028 228467 202078 228977
rect 202398 228467 204448 228977
rect 205028 228467 206851 228977
rect 218272 227877 220172 228367
rect 220752 227877 222802 228367
rect 223122 227877 225172 228367
rect 225828 227877 227878 228367
rect 228198 227877 230248 228367
rect 230828 227877 232655 228367
rect 192472 227255 194372 227765
rect 194952 227255 197002 227765
rect 197322 227255 199372 227765
rect 200028 227255 202078 227765
rect 202398 227255 204448 227765
rect 205028 227255 206851 227765
rect 218272 226665 220172 227155
rect 220752 226665 222802 227155
rect 223122 226665 225172 227155
rect 225828 226665 227878 227155
rect 228198 226665 230248 227155
rect 230828 226665 232655 227155
rect 192472 226043 194372 226553
rect 194952 226043 197002 226553
rect 197322 226043 199372 226553
rect 200028 226043 202078 226553
rect 202398 226043 204448 226553
rect 205028 226043 206851 226553
rect 218272 225453 220172 225943
rect 220752 225453 222802 225943
rect 223122 225453 225172 225943
rect 225828 225453 227878 225943
rect 228198 225453 230248 225943
rect 230828 225453 232655 225943
rect 192472 224831 194372 225341
rect 194952 224831 197002 225341
rect 197322 224831 199372 225341
rect 200028 224831 202078 225341
rect 202398 224831 204448 225341
rect 205028 224831 206851 225341
rect 218272 224241 220172 224731
rect 220752 224241 222802 224731
rect 223122 224241 225172 224731
rect 225828 224241 227878 224731
rect 228198 224241 230248 224731
rect 230828 224241 232655 224731
rect 192472 223619 194372 224129
rect 194952 223619 197002 224129
rect 197322 223619 199372 224129
rect 200028 223619 202078 224129
rect 202398 223619 204448 224129
rect 205028 223619 206851 224129
rect 218272 223029 220172 223519
rect 220752 223029 222802 223519
rect 223122 223029 225172 223519
rect 225828 223029 227878 223519
rect 228198 223029 230248 223519
rect 230828 223029 232655 223519
rect 192472 222407 194372 222917
rect 194952 222407 197002 222917
rect 197322 222407 199372 222917
rect 200028 222407 202078 222917
rect 202398 222407 204448 222917
rect 205028 222407 206851 222917
rect 218272 221817 220172 222307
rect 220752 221817 222802 222307
rect 223122 221817 225172 222307
rect 225828 221817 227878 222307
rect 228198 221817 230248 222307
rect 230828 221817 232655 222307
rect 192472 221195 194372 221705
rect 194952 221195 197002 221705
rect 197322 221195 199372 221705
rect 200028 221195 202078 221705
rect 202398 221195 204448 221705
rect 205028 221195 206851 221705
rect 218272 220605 220172 221095
rect 220752 220605 222802 221095
rect 223122 220605 225172 221095
rect 225828 220605 227878 221095
rect 228198 220605 230248 221095
rect 230828 220605 232655 221095
rect 192472 219983 194372 220493
rect 194952 219983 197002 220493
rect 197322 219983 199372 220493
rect 200028 219983 202078 220493
rect 202398 219983 204448 220493
rect 205028 219983 206851 220493
rect 218272 219393 220172 219883
rect 220752 219393 222802 219883
rect 223122 219393 225172 219883
rect 225828 219393 227878 219883
rect 228198 219393 230248 219883
rect 230828 219393 232655 219883
rect 192472 218771 194372 219281
rect 194952 218771 197002 219281
rect 197322 218771 199372 219281
rect 200028 218771 202078 219281
rect 202398 218771 204448 219281
rect 205028 218771 206851 219281
rect 218272 218181 220172 218671
rect 220752 218181 222802 218671
rect 223122 218181 225172 218671
rect 225828 218181 227878 218671
rect 228198 218181 230248 218671
rect 230828 218181 232655 218671
rect 192472 217559 194372 218069
rect 194952 217559 197002 218069
rect 197322 217559 199372 218069
rect 200028 217559 202078 218069
rect 202398 217559 204448 218069
rect 205028 217559 206851 218069
rect 75272 217039 75332 217098
rect 218272 216969 220172 217459
rect 220752 216969 222802 217459
rect 223122 216969 225172 217459
rect 225828 216969 227878 217459
rect 228198 216969 230248 217459
rect 230828 216969 232655 217459
rect 192472 216347 194372 216857
rect 194952 216347 197002 216857
rect 197322 216347 199372 216857
rect 200028 216347 202078 216857
rect 202398 216347 204448 216857
rect 205028 216347 206851 216857
rect 75392 216166 75452 216225
rect 218272 215757 220172 216247
rect 220752 215757 222802 216247
rect 223122 215757 225172 216247
rect 225828 215757 227878 216247
rect 228198 215757 230248 216247
rect 230828 215757 232655 216247
rect 192472 215135 194372 215645
rect 194952 215135 197002 215645
rect 197322 215135 199372 215645
rect 200028 215135 202078 215645
rect 202398 215135 204448 215645
rect 205028 215135 206851 215645
rect 218272 214545 220172 215035
rect 220752 214545 222802 215035
rect 223122 214545 225172 215035
rect 225828 214545 227878 215035
rect 228198 214545 230248 215035
rect 230828 214545 232655 215035
rect 192472 213923 194372 214433
rect 194952 213923 197002 214433
rect 197322 213923 199372 214433
rect 200028 213923 202078 214433
rect 202398 213923 204448 214433
rect 205028 213923 206851 214433
rect 218272 213333 220172 213823
rect 220752 213333 222802 213823
rect 223122 213333 225172 213823
rect 225828 213333 227878 213823
rect 228198 213333 230248 213823
rect 230828 213333 232655 213823
rect 192472 212711 194372 213221
rect 194952 212711 197002 213221
rect 197322 212711 199372 213221
rect 200028 212711 202078 213221
rect 202398 212711 204448 213221
rect 205028 212711 206851 213221
rect 218272 212121 220172 212611
rect 220752 212121 222802 212611
rect 223122 212121 225172 212611
rect 225828 212121 227878 212611
rect 228198 212121 230248 212611
rect 230828 212121 232655 212611
rect 192472 211499 194372 212009
rect 194952 211499 197002 212009
rect 197322 211499 199372 212009
rect 200028 211499 202078 212009
rect 202398 211499 204448 212009
rect 205028 211499 206851 212009
rect 218272 210876 220172 211576
rect 220752 210876 222802 211576
rect 223122 210876 225172 211576
rect 225828 210876 227878 211576
rect 228198 210876 230248 211576
rect 230828 210876 232655 211576
rect 192472 210287 194372 210797
rect 194952 210287 197002 210797
rect 197322 210287 199372 210797
rect 200028 210287 202078 210797
rect 202398 210287 204448 210797
rect 205028 210287 206851 210797
rect 218272 209697 220172 210187
rect 220752 209697 222802 210187
rect 223122 209697 225172 210187
rect 225828 209697 227878 210187
rect 228198 209697 230248 210187
rect 230828 209697 232655 210187
rect 192472 209095 194372 209585
rect 194952 209095 197002 209585
rect 197322 209095 199372 209585
rect 200028 209095 202078 209585
rect 202398 209095 204448 209585
rect 205028 209095 206851 209585
rect 218272 208485 220172 208975
rect 220752 208485 222802 208975
rect 223122 208485 225172 208975
rect 225828 208485 227878 208975
rect 228198 208485 230248 208975
rect 230828 208485 232655 208975
rect 192472 207883 194372 208373
rect 194952 207883 197002 208373
rect 197322 207883 199372 208373
rect 200028 207883 202078 208373
rect 202398 207883 204448 208373
rect 205028 207883 206851 208373
rect 218272 207273 220172 207763
rect 220752 207273 222802 207763
rect 223122 207273 225172 207763
rect 225828 207273 227878 207763
rect 228198 207273 230248 207763
rect 230828 207273 232655 207763
rect 192472 206671 194372 207161
rect 194952 206671 197002 207161
rect 197322 206671 199372 207161
rect 200028 206671 202078 207161
rect 202398 206671 204448 207161
rect 205028 206671 206851 207161
rect 218272 206061 220172 206551
rect 220752 206061 222802 206551
rect 223122 206061 225172 206551
rect 225828 206061 227878 206551
rect 228198 206061 230248 206551
rect 230828 206061 232655 206551
rect 192472 205459 194372 205949
rect 194952 205459 197002 205949
rect 197322 205459 199372 205949
rect 200028 205459 202078 205949
rect 202398 205459 204448 205949
rect 205028 205459 206851 205949
rect 218272 204849 220172 205339
rect 220752 204849 222802 205339
rect 223122 204849 225172 205339
rect 225828 204849 227878 205339
rect 228198 204849 230248 205339
rect 230828 204849 232655 205339
rect 192472 204247 194372 204737
rect 194952 204247 197002 204737
rect 197322 204247 199372 204737
rect 200028 204247 202078 204737
rect 202398 204247 204448 204737
rect 205028 204247 206851 204737
rect 218272 203637 220172 204127
rect 220752 203637 222802 204127
rect 223122 203637 225172 204127
rect 225828 203637 227878 204127
rect 228198 203637 230248 204127
rect 230828 203637 232655 204127
rect 192472 203035 194372 203525
rect 194952 203035 197002 203525
rect 197322 203035 199372 203525
rect 200028 203035 202078 203525
rect 202398 203035 204448 203525
rect 205028 203035 206851 203525
rect 218272 202425 220172 202915
rect 220752 202425 222802 202915
rect 223122 202425 225172 202915
rect 225828 202425 227878 202915
rect 228198 202425 230248 202915
rect 230828 202425 232655 202915
rect 192472 201823 194372 202313
rect 194952 201823 197002 202313
rect 197322 201823 199372 202313
rect 200028 201823 202078 202313
rect 202398 201823 204448 202313
rect 205028 201823 206851 202313
rect 218272 201213 220172 201703
rect 220752 201213 222802 201703
rect 223122 201213 225172 201703
rect 225828 201213 227878 201703
rect 228198 201213 230248 201703
rect 230828 201213 232655 201703
rect 192472 200611 194372 201101
rect 194952 200611 197002 201101
rect 197322 200611 199372 201101
rect 200028 200611 202078 201101
rect 202398 200611 204448 201101
rect 205028 200611 206851 201101
rect 218272 200001 220172 200491
rect 220752 200001 222802 200491
rect 223122 200001 225172 200491
rect 225828 200001 227878 200491
rect 228198 200001 230248 200491
rect 230828 200001 232655 200491
rect 192472 199399 194372 199889
rect 194952 199399 197002 199889
rect 197322 199399 199372 199889
rect 200028 199399 202078 199889
rect 202398 199399 204448 199889
rect 205028 199399 206851 199889
rect 218272 198789 220172 199279
rect 220752 198789 222802 199279
rect 223122 198789 225172 199279
rect 225828 198789 227878 199279
rect 228198 198789 230248 199279
rect 230828 198789 232655 199279
rect 192472 198187 194372 198677
rect 194952 198187 197002 198677
rect 197322 198187 199372 198677
rect 200028 198187 202078 198677
rect 202398 198187 204448 198677
rect 205028 198187 206851 198677
rect 218272 197577 220172 198067
rect 220752 197577 222802 198067
rect 223122 197577 225172 198067
rect 225828 197577 227878 198067
rect 228198 197577 230248 198067
rect 230828 197577 232655 198067
rect 192472 196975 194372 197465
rect 194952 196975 197002 197465
rect 197322 196975 199372 197465
rect 200028 196975 202078 197465
rect 202398 196975 204448 197465
rect 205028 196975 206851 197465
rect 218272 196365 220172 196855
rect 220752 196365 222802 196855
rect 223122 196365 225172 196855
rect 225828 196365 227878 196855
rect 228198 196365 230248 196855
rect 230828 196365 232655 196855
rect 192472 195763 194372 196253
rect 194952 195763 197002 196253
rect 197322 195763 199372 196253
rect 200028 195763 202078 196253
rect 202398 195763 204448 196253
rect 205028 195763 206851 196253
rect 218272 195153 220172 195643
rect 220752 195153 222802 195643
rect 223122 195153 225172 195643
rect 225828 195153 227878 195643
rect 228198 195153 230248 195643
rect 230828 195153 232655 195643
rect 192472 194551 194372 195041
rect 194952 194551 197002 195041
rect 197322 194551 199372 195041
rect 200028 194551 202078 195041
rect 202398 194551 204448 195041
rect 205028 194551 206851 195041
rect 218272 193941 220172 194431
rect 220752 193941 222802 194431
rect 223122 193941 225172 194431
rect 225828 193941 227878 194431
rect 228198 193941 230248 194431
rect 230828 193941 232655 194431
rect 192472 193339 194372 193829
rect 194952 193339 197002 193829
rect 197322 193339 199372 193829
rect 200028 193339 202078 193829
rect 202398 193339 204448 193829
rect 205028 193339 206851 193829
rect 218272 192729 220172 193219
rect 220752 192729 222802 193219
rect 223122 192729 225172 193219
rect 225828 192729 227878 193219
rect 228198 192729 230248 193219
rect 230828 192729 232655 193219
rect 192472 192127 194372 192617
rect 194952 192127 197002 192617
rect 197322 192127 199372 192617
rect 200028 192127 202078 192617
rect 202398 192127 204448 192617
rect 205028 192127 206851 192617
rect 218272 191517 220172 192007
rect 220752 191517 222802 192007
rect 223122 191517 225172 192007
rect 225828 191517 227878 192007
rect 228198 191517 230248 192007
rect 230828 191517 232655 192007
rect 192472 190915 194372 191405
rect 194952 190915 197002 191405
rect 197322 190915 199372 191405
rect 200028 190915 202078 191405
rect 202398 190915 204448 191405
rect 205028 190915 206851 191405
rect 579472 190983 581372 191683
rect 581952 190983 584002 191683
rect 584322 190983 586372 191683
rect 587028 190983 589078 191683
rect 589398 190983 591448 191683
rect 592028 190983 593928 191683
rect 218272 190305 220172 190795
rect 220752 190305 222802 190795
rect 223122 190305 225172 190795
rect 225828 190305 227878 190795
rect 228198 190305 230248 190795
rect 230828 190305 232655 190795
rect 553672 190394 555572 190904
rect 556152 190394 558202 190904
rect 558522 190394 560572 190904
rect 561228 190394 563278 190904
rect 563598 190394 565648 190904
rect 566228 190394 568128 190904
rect 192472 189703 194372 190193
rect 194952 189703 197002 190193
rect 197322 189703 199372 190193
rect 200028 189703 202078 190193
rect 202398 189703 204448 190193
rect 205028 189703 206851 190193
rect 579472 189804 581372 190294
rect 581952 189804 584002 190294
rect 584322 189804 586372 190294
rect 587028 189804 589078 190294
rect 589398 189804 591448 190294
rect 592028 189804 593928 190294
rect 218272 189093 220172 189583
rect 220752 189093 222802 189583
rect 223122 189093 225172 189583
rect 225828 189093 227878 189583
rect 228198 189093 230248 189583
rect 230828 189093 232655 189583
rect 553672 189202 555572 189692
rect 556152 189202 558202 189692
rect 558522 189202 560572 189692
rect 561228 189202 563278 189692
rect 563598 189202 565648 189692
rect 566228 189202 568128 189692
rect 75272 188839 75332 188898
rect 192472 188491 194372 188981
rect 194952 188491 197002 188981
rect 197322 188491 199372 188981
rect 200028 188491 202078 188981
rect 202398 188491 204448 188981
rect 205028 188491 206851 188981
rect 579472 188592 581372 189082
rect 581952 188592 584002 189082
rect 584322 188592 586372 189082
rect 587028 188592 589078 189082
rect 589398 188592 591448 189082
rect 592028 188592 593928 189082
rect 75272 187966 75332 188025
rect 218272 187881 220172 188371
rect 220752 187881 222802 188371
rect 223122 187881 225172 188371
rect 225828 187881 227878 188371
rect 228198 187881 230248 188371
rect 230828 187881 232655 188371
rect 553672 187990 555572 188480
rect 556152 187990 558202 188480
rect 558522 187990 560572 188480
rect 561228 187990 563278 188480
rect 563598 187990 565648 188480
rect 566228 187990 568128 188480
rect 192472 187279 194372 187769
rect 194952 187279 197002 187769
rect 197322 187279 199372 187769
rect 200028 187279 202078 187769
rect 202398 187279 204448 187769
rect 205028 187279 206851 187769
rect 579472 187380 581372 187870
rect 581952 187380 584002 187870
rect 584322 187380 586372 187870
rect 587028 187380 589078 187870
rect 589398 187380 591448 187870
rect 592028 187380 593928 187870
rect 218272 186669 220172 187159
rect 220752 186669 222802 187159
rect 223122 186669 225172 187159
rect 225828 186669 227878 187159
rect 228198 186669 230248 187159
rect 230828 186669 232655 187159
rect 553672 186778 555572 187268
rect 556152 186778 558202 187268
rect 558522 186778 560572 187268
rect 561228 186778 563278 187268
rect 563598 186778 565648 187268
rect 566228 186778 568128 187268
rect 192472 186067 194372 186557
rect 194952 186067 197002 186557
rect 197322 186067 199372 186557
rect 200028 186067 202078 186557
rect 202398 186067 204448 186557
rect 205028 186067 206851 186557
rect 579472 186168 581372 186658
rect 581952 186168 584002 186658
rect 584322 186168 586372 186658
rect 587028 186168 589078 186658
rect 589398 186168 591448 186658
rect 592028 186168 593928 186658
rect 218272 185457 220172 185947
rect 220752 185457 222802 185947
rect 223122 185457 225172 185947
rect 225828 185457 227878 185947
rect 228198 185457 230248 185947
rect 230828 185457 232655 185947
rect 553672 185566 555572 186056
rect 556152 185566 558202 186056
rect 558522 185566 560572 186056
rect 561228 185566 563278 186056
rect 563598 185566 565648 186056
rect 566228 185566 568128 186056
rect 192472 184855 194372 185345
rect 194952 184855 197002 185345
rect 197322 184855 199372 185345
rect 200028 184855 202078 185345
rect 202398 184855 204448 185345
rect 205028 184855 206851 185345
rect 579472 184956 581372 185446
rect 581952 184956 584002 185446
rect 584322 184956 586372 185446
rect 587028 184956 589078 185446
rect 589398 184956 591448 185446
rect 592028 184956 593928 185446
rect 218272 184245 220172 184735
rect 220752 184245 222802 184735
rect 223122 184245 225172 184735
rect 225828 184245 227878 184735
rect 228198 184245 230248 184735
rect 230828 184245 232655 184735
rect 553672 184354 555572 184844
rect 556152 184354 558202 184844
rect 558522 184354 560572 184844
rect 561228 184354 563278 184844
rect 563598 184354 565648 184844
rect 566228 184354 568128 184844
rect 192472 183643 194372 184133
rect 194952 183643 197002 184133
rect 197322 183643 199372 184133
rect 200028 183643 202078 184133
rect 202398 183643 204448 184133
rect 205028 183643 206851 184133
rect 579472 183744 581372 184234
rect 581952 183744 584002 184234
rect 584322 183744 586372 184234
rect 587028 183744 589078 184234
rect 589398 183744 591448 184234
rect 592028 183744 593928 184234
rect 218272 183033 220172 183523
rect 220752 183033 222802 183523
rect 223122 183033 225172 183523
rect 225828 183033 227878 183523
rect 228198 183033 230248 183523
rect 230828 183033 232655 183523
rect 553672 183142 555572 183632
rect 556152 183142 558202 183632
rect 558522 183142 560572 183632
rect 561228 183142 563278 183632
rect 563598 183142 565648 183632
rect 566228 183142 568128 183632
rect 192472 182431 194372 182921
rect 194952 182431 197002 182921
rect 197322 182431 199372 182921
rect 200028 182431 202078 182921
rect 202398 182431 204448 182921
rect 205028 182431 206851 182921
rect 579472 182532 581372 183022
rect 581952 182532 584002 183022
rect 584322 182532 586372 183022
rect 587028 182532 589078 183022
rect 589398 182532 591448 183022
rect 592028 182532 593928 183022
rect 218272 181821 220172 182311
rect 220752 181821 222802 182311
rect 223122 181821 225172 182311
rect 225828 181821 227878 182311
rect 228198 181821 230248 182311
rect 230828 181821 232655 182311
rect 553672 181930 555572 182420
rect 556152 181930 558202 182420
rect 558522 181930 560572 182420
rect 561228 181930 563278 182420
rect 563598 181930 565648 182420
rect 566228 181930 568128 182420
rect 192472 181219 194372 181709
rect 194952 181219 197002 181709
rect 197322 181219 199372 181709
rect 200028 181219 202078 181709
rect 202398 181219 204448 181709
rect 205028 181219 206851 181709
rect 579472 181320 581372 181810
rect 581952 181320 584002 181810
rect 584322 181320 586372 181810
rect 587028 181320 589078 181810
rect 589398 181320 591448 181810
rect 592028 181320 593928 181810
rect 218272 180609 220172 181099
rect 220752 180609 222802 181099
rect 223122 180609 225172 181099
rect 225828 180609 227878 181099
rect 228198 180609 230248 181099
rect 230828 180609 232655 181099
rect 553672 180718 555572 181208
rect 556152 180718 558202 181208
rect 558522 180718 560572 181208
rect 561228 180718 563278 181208
rect 563598 180718 565648 181208
rect 566228 180718 568128 181208
rect 192472 180007 194372 180497
rect 194952 180007 197002 180497
rect 197322 180007 199372 180497
rect 200028 180007 202078 180497
rect 202398 180007 204448 180497
rect 205028 180007 206851 180497
rect 579472 180108 581372 180598
rect 581952 180108 584002 180598
rect 584322 180108 586372 180598
rect 587028 180108 589078 180598
rect 589398 180108 591448 180598
rect 592028 180108 593928 180598
rect 218272 179397 220172 179887
rect 220752 179397 222802 179887
rect 223122 179397 225172 179887
rect 225828 179397 227878 179887
rect 228198 179397 230248 179887
rect 230828 179397 232655 179887
rect 553672 179506 555572 179996
rect 556152 179506 558202 179996
rect 558522 179506 560572 179996
rect 561228 179506 563278 179996
rect 563598 179506 565648 179996
rect 566228 179506 568128 179996
rect 192472 178795 194372 179285
rect 194952 178795 197002 179285
rect 197322 178795 199372 179285
rect 200028 178795 202078 179285
rect 202398 178795 204448 179285
rect 205028 178795 206851 179285
rect 579472 178896 581372 179386
rect 581952 178896 584002 179386
rect 584322 178896 586372 179386
rect 587028 178896 589078 179386
rect 589398 178896 591448 179386
rect 592028 178896 593928 179386
rect 218272 178185 220172 178675
rect 220752 178185 222802 178675
rect 223122 178185 225172 178675
rect 225828 178185 227878 178675
rect 228198 178185 230248 178675
rect 230828 178185 232655 178675
rect 553672 178294 555572 178784
rect 556152 178294 558202 178784
rect 558522 178294 560572 178784
rect 561228 178294 563278 178784
rect 563598 178294 565648 178784
rect 566228 178294 568128 178784
rect 192472 177583 194372 178073
rect 194952 177583 197002 178073
rect 197322 177583 199372 178073
rect 200028 177583 202078 178073
rect 202398 177583 204448 178073
rect 205028 177583 206851 178073
rect 579472 177684 581372 178174
rect 581952 177684 584002 178174
rect 584322 177684 586372 178174
rect 587028 177684 589078 178174
rect 589398 177684 591448 178174
rect 592028 177684 593928 178174
rect 218272 176973 220172 177463
rect 220752 176973 222802 177463
rect 223122 176973 225172 177463
rect 225828 176973 227878 177463
rect 228198 176973 230248 177463
rect 230828 176973 232655 177463
rect 553672 177082 555572 177572
rect 556152 177082 558202 177572
rect 558522 177082 560572 177572
rect 561228 177082 563278 177572
rect 563598 177082 565648 177572
rect 566228 177082 568128 177572
rect 192472 176371 194372 176861
rect 194952 176371 197002 176861
rect 197322 176371 199372 176861
rect 200028 176371 202078 176861
rect 202398 176371 204448 176861
rect 205028 176371 206851 176861
rect 579472 176472 581372 176962
rect 581952 176472 584002 176962
rect 584322 176472 586372 176962
rect 587028 176472 589078 176962
rect 589398 176472 591448 176962
rect 592028 176472 593928 176962
rect 218272 175761 220172 176251
rect 220752 175761 222802 176251
rect 223122 175761 225172 176251
rect 225828 175761 227878 176251
rect 228198 175761 230248 176251
rect 230828 175761 232655 176251
rect 553672 175870 555572 176360
rect 556152 175870 558202 176360
rect 558522 175870 560572 176360
rect 561228 175870 563278 176360
rect 563598 175870 565648 176360
rect 566228 175870 568128 176360
rect 192472 175159 194372 175649
rect 194952 175159 197002 175649
rect 197322 175159 199372 175649
rect 200028 175159 202078 175649
rect 202398 175159 204448 175649
rect 205028 175159 206851 175649
rect 579472 175260 581372 175750
rect 581952 175260 584002 175750
rect 584322 175260 586372 175750
rect 587028 175260 589078 175750
rect 589398 175260 591448 175750
rect 592028 175260 593928 175750
rect 218272 174549 220172 175039
rect 220752 174549 222802 175039
rect 223122 174549 225172 175039
rect 225828 174549 227878 175039
rect 228198 174549 230248 175039
rect 230828 174549 232655 175039
rect 553672 174658 555572 175148
rect 556152 174658 558202 175148
rect 558522 174658 560572 175148
rect 561228 174658 563278 175148
rect 563598 174658 565648 175148
rect 566228 174658 568128 175148
rect 192472 173947 194372 174437
rect 194952 173947 197002 174437
rect 197322 173947 199372 174437
rect 200028 173947 202078 174437
rect 202398 173947 204448 174437
rect 205028 173947 206851 174437
rect 579472 174048 581372 174538
rect 581952 174048 584002 174538
rect 584322 174048 586372 174538
rect 587028 174048 589078 174538
rect 589398 174048 591448 174538
rect 592028 174048 593928 174538
rect 218272 173337 220172 173827
rect 220752 173337 222802 173827
rect 223122 173337 225172 173827
rect 225828 173337 227878 173827
rect 228198 173337 230248 173827
rect 230828 173337 232655 173827
rect 553672 173446 555572 173936
rect 556152 173446 558202 173936
rect 558522 173446 560572 173936
rect 561228 173446 563278 173936
rect 563598 173446 565648 173936
rect 566228 173446 568128 173936
rect 192472 172735 194372 173225
rect 194952 172735 197002 173225
rect 197322 172735 199372 173225
rect 200028 172735 202078 173225
rect 202398 172735 204448 173225
rect 205028 172735 206851 173225
rect 579472 172836 581372 173326
rect 581952 172836 584002 173326
rect 584322 172836 586372 173326
rect 587028 172836 589078 173326
rect 589398 172836 591448 173326
rect 592028 172836 593928 173326
rect 218272 172125 220172 172615
rect 220752 172125 222802 172615
rect 223122 172125 225172 172615
rect 225828 172125 227878 172615
rect 228198 172125 230248 172615
rect 230828 172125 232655 172615
rect 553672 172234 555572 172724
rect 556152 172234 558202 172724
rect 558522 172234 560572 172724
rect 561228 172234 563278 172724
rect 563598 172234 565648 172724
rect 566228 172234 568128 172724
rect 192472 171523 194372 172013
rect 194952 171523 197002 172013
rect 197322 171523 199372 172013
rect 200028 171523 202078 172013
rect 202398 171523 204448 172013
rect 205028 171523 206851 172013
rect 579472 171624 581372 172114
rect 581952 171624 584002 172114
rect 584322 171624 586372 172114
rect 587028 171624 589078 172114
rect 589398 171624 591448 172114
rect 592028 171624 593928 172114
rect 218272 170913 220172 171403
rect 220752 170913 222802 171403
rect 223122 170913 225172 171403
rect 225828 170913 227878 171403
rect 228198 170913 230248 171403
rect 230828 170913 232655 171403
rect 553672 171022 555572 171512
rect 556152 171022 558202 171512
rect 558522 171022 560572 171512
rect 561228 171022 563278 171512
rect 563598 171022 565648 171512
rect 566228 171022 568128 171512
rect 192472 170027 194372 170630
rect 194952 170027 197002 170630
rect 197322 170027 199372 170630
rect 200028 170027 202078 170630
rect 202398 170027 204448 170630
rect 205028 170027 206851 170630
rect 579472 170412 581372 170902
rect 581952 170412 584002 170902
rect 584322 170412 586372 170902
rect 587028 170412 589078 170902
rect 589398 170412 591448 170902
rect 592028 170412 593928 170902
rect 218272 166792 220172 169740
rect 220752 166792 222802 169740
rect 223122 166792 225172 169740
rect 225828 166792 227878 169740
rect 228198 166792 230248 169740
rect 230828 166792 232655 169740
rect 553672 169526 555572 170129
rect 556152 169526 558202 170129
rect 558522 169526 560572 170129
rect 561228 169526 563278 170129
rect 563598 169526 565648 170129
rect 566228 169526 568128 170129
rect 192472 165136 194372 166524
rect 194952 165136 197002 166524
rect 197322 165136 199372 166524
rect 200028 165136 202078 166524
rect 202398 165136 204448 166524
rect 205028 165136 206851 166524
rect 579472 166291 581372 169239
rect 581952 166291 584002 169239
rect 584322 166291 586372 169239
rect 587028 166291 589078 169239
rect 589398 166291 591448 169239
rect 592028 166291 593928 169239
rect 553672 164635 555572 166023
rect 556152 164635 558202 166023
rect 558522 164635 560572 166023
rect 561228 164635 563278 166023
rect 563598 164635 565648 166023
rect 566228 164635 568128 166023
rect 218272 162728 220172 163429
rect 220752 162728 222802 163429
rect 223122 162728 225172 163429
rect 225828 162728 227878 163429
rect 228198 162728 230248 163429
rect 230828 162728 232655 163429
rect 192472 161629 194372 162330
rect 194952 161629 197002 162330
rect 197322 161629 199372 162330
rect 200028 161629 202078 162330
rect 202398 161629 204448 162330
rect 205028 161629 206851 162330
rect 579472 162227 581372 162928
rect 581952 162227 584002 162928
rect 584322 162227 586372 162928
rect 587028 162227 589078 162928
rect 589398 162227 591448 162928
rect 592028 162227 593928 162928
rect 75272 160639 75332 160698
rect 75272 159766 75332 159825
rect 218272 159399 220172 161308
rect 220752 159399 222802 161308
rect 223122 159399 225172 161308
rect 225828 159399 227878 161308
rect 228198 159399 230248 161308
rect 230828 159399 232655 161308
rect 553672 161128 555572 161829
rect 556152 161128 558202 161829
rect 558522 161128 560572 161829
rect 561228 161128 563278 161829
rect 563598 161128 565648 161829
rect 566228 161128 568128 161829
rect 192472 157348 194372 159200
rect 194952 157348 197002 159200
rect 197322 157348 199372 159200
rect 200028 157348 202078 159200
rect 202398 157348 204448 159200
rect 205028 157348 206851 159200
rect 579472 158898 581372 160807
rect 581952 158898 584002 160807
rect 584322 158898 586372 160807
rect 587028 158898 589078 160807
rect 589398 158898 591448 160807
rect 592028 158898 593928 160807
rect 218272 155760 220172 157222
rect 220752 155760 222802 157222
rect 223122 155760 225172 157222
rect 225828 155760 227878 157222
rect 228198 155760 230248 157222
rect 230828 155760 232655 157222
rect 553672 156847 555572 158699
rect 556152 156847 558202 158699
rect 558522 156847 560572 158699
rect 561228 156847 563278 158699
rect 563598 156847 565648 158699
rect 566228 156847 568128 158699
rect 192472 154481 194372 155404
rect 194952 154481 197002 155404
rect 197322 154481 199372 155404
rect 200028 154481 202078 155404
rect 202398 154481 204448 155404
rect 205028 154481 206851 155404
rect 579472 155259 581372 156721
rect 581952 155259 584002 156721
rect 584322 155259 586372 156721
rect 587028 155259 589078 156721
rect 589398 155259 591448 156721
rect 592028 155259 593928 156721
rect 218272 153063 220172 154018
rect 220752 153063 222802 154018
rect 223122 153063 225172 154018
rect 225828 153063 227878 154018
rect 228198 153063 230248 154018
rect 230828 153063 232655 154018
rect 553672 153980 555572 154903
rect 556152 153980 558202 154903
rect 558522 153980 560572 154903
rect 561228 153980 563278 154903
rect 563598 153980 565648 154903
rect 566228 153980 568128 154903
rect 192472 151720 194372 152851
rect 194952 151720 197002 152851
rect 197322 151720 199372 152851
rect 200028 151720 202078 152851
rect 202398 151720 204448 152851
rect 205028 151720 206851 152851
rect 579472 152562 581372 153517
rect 581952 152562 584002 153517
rect 584322 152562 586372 153517
rect 587028 152562 589078 153517
rect 589398 152562 591448 153517
rect 592028 152562 593928 153517
rect 218272 150599 220172 151628
rect 220752 150599 222802 151628
rect 223122 150599 225172 151628
rect 225828 150599 227878 151628
rect 228198 150599 230248 151628
rect 230828 150599 232655 151628
rect 553672 151219 555572 152350
rect 556152 151219 558202 152350
rect 558522 151219 560572 152350
rect 561228 151219 563278 152350
rect 563598 151219 565648 152350
rect 566228 151219 568128 152350
rect 192472 149508 194372 150397
rect 194952 149508 197002 150397
rect 197322 149508 199372 150397
rect 200028 149508 202078 150397
rect 202398 149508 204448 150397
rect 205028 149508 206851 150397
rect 459446 150035 460246 150332
rect 579472 150098 581372 151127
rect 581952 150098 584002 151127
rect 584322 150098 586372 151127
rect 587028 150098 589078 151127
rect 589398 150098 591448 151127
rect 592028 150098 593928 151127
rect 328649 149896 329463 150030
rect 460979 149414 461779 149711
rect 218272 148620 220172 149320
rect 220752 148620 222802 149320
rect 223122 148620 225172 149320
rect 225828 148620 227878 149320
rect 228198 148620 230248 149320
rect 230828 148620 232655 149320
rect 327021 149098 327835 149232
rect 553672 149007 555572 149896
rect 556152 149007 558202 149896
rect 558522 149007 560572 149896
rect 561228 149007 563278 149896
rect 563598 149007 565648 149896
rect 566228 149007 568128 149896
rect 579472 148119 581372 148819
rect 581952 148119 584002 148819
rect 584322 148119 586372 148819
rect 587028 148119 589078 148819
rect 589398 148119 591448 148819
rect 592028 148119 593928 148819
rect 218272 86550 220172 87078
<< metal4 >>
rect 218272 415428 220172 417503
rect 218272 412948 220172 413528
rect 218272 410578 220172 410898
rect 218272 407872 220172 408528
rect 218272 405502 220172 405822
rect 218272 402872 220172 403452
rect 192472 387228 194372 390292
rect 192472 384748 194372 385328
rect 192472 382378 194372 382698
rect 192472 379672 194372 380328
rect 192472 377302 194372 377622
rect 192472 374672 194372 375252
rect 192472 249581 194372 372772
rect 192472 248369 194372 249071
rect 192472 247157 194372 247859
rect 192472 245945 194372 246647
rect 192472 244733 194372 245435
rect 192472 243521 194372 244223
rect 192472 242309 194372 243011
rect 192472 241097 194372 241799
rect 192472 239885 194372 240587
rect 192472 238673 194372 239375
rect 192472 237461 194372 238163
rect 192472 236249 194372 236951
rect 192472 235037 194372 235739
rect 192472 233825 194372 234527
rect 192472 232613 194372 233315
rect 192472 231401 194372 232103
rect 192472 230189 194372 230891
rect 192472 228977 194372 229679
rect 192472 227765 194372 228467
rect 192472 226553 194372 227255
rect 192472 225341 194372 226043
rect 192472 224129 194372 224831
rect 192472 222917 194372 223619
rect 192472 221705 194372 222407
rect 192472 220493 194372 221195
rect 192472 219281 194372 219983
rect 192472 218069 194372 218771
rect 192472 216857 194372 217559
rect 192472 215645 194372 216347
rect 192472 214433 194372 215135
rect 192472 213221 194372 213923
rect 192472 212009 194372 212711
rect 192472 210797 194372 211499
rect 192472 209585 194372 210287
rect 192472 208373 194372 209095
rect 192472 207161 194372 207883
rect 192472 205949 194372 206671
rect 192472 204737 194372 205459
rect 192472 203525 194372 204247
rect 192472 202313 194372 203035
rect 192472 201101 194372 201823
rect 192472 199889 194372 200611
rect 192472 198677 194372 199399
rect 192472 197465 194372 198187
rect 192472 196253 194372 196975
rect 192472 195041 194372 195763
rect 192472 193829 194372 194551
rect 192472 192617 194372 193339
rect 192472 191405 194372 192127
rect 192472 190193 194372 190915
rect 192472 188981 194372 189703
rect 192472 187769 194372 188491
rect 192472 186557 194372 187279
rect 192472 185345 194372 186067
rect 192472 184133 194372 184855
rect 192472 182921 194372 183643
rect 192472 181709 194372 182431
rect 192472 180497 194372 181219
rect 192472 179285 194372 180007
rect 192472 178073 194372 178795
rect 192472 176861 194372 177583
rect 192472 175649 194372 176371
rect 192472 174437 194372 175159
rect 192472 173225 194372 173947
rect 192472 172013 194372 172735
rect 192472 170630 194372 171523
rect 192472 166524 194372 170027
rect 192472 162330 194372 165136
rect 192472 159200 194372 161629
rect 192472 155404 194372 157348
rect 192472 152851 194372 154481
rect 192472 150397 194372 151720
rect 192472 105228 194372 149508
rect 192472 102748 194372 103328
rect 192472 100378 194372 100698
rect 192472 97672 194372 98328
rect 192472 95302 194372 95622
rect 192472 92672 194372 93252
rect 192472 75400 194372 90772
rect 194952 387228 197002 390292
rect 194952 384748 197002 385328
rect 194952 382378 197002 382698
rect 194952 379672 197002 380328
rect 194952 377302 197002 377622
rect 194952 374672 197002 375252
rect 194952 249581 197002 372772
rect 194952 248369 197002 249071
rect 194952 247157 197002 247859
rect 194952 245945 197002 246647
rect 194952 244733 197002 245435
rect 194952 243521 197002 244223
rect 194952 242309 197002 243011
rect 194952 241097 197002 241799
rect 194952 239885 197002 240587
rect 194952 238673 197002 239375
rect 194952 237461 197002 238163
rect 194952 236249 197002 236951
rect 194952 235037 197002 235739
rect 194952 233825 197002 234527
rect 194952 232613 197002 233315
rect 194952 231401 197002 232103
rect 194952 230189 197002 230891
rect 194952 228977 197002 229679
rect 194952 227765 197002 228467
rect 194952 226553 197002 227255
rect 194952 225341 197002 226043
rect 194952 224129 197002 224831
rect 194952 222917 197002 223619
rect 194952 221705 197002 222407
rect 194952 220493 197002 221195
rect 194952 219281 197002 219983
rect 194952 218069 197002 218771
rect 194952 216857 197002 217559
rect 194952 215645 197002 216347
rect 194952 214433 197002 215135
rect 194952 213221 197002 213923
rect 194952 212009 197002 212711
rect 194952 210797 197002 211499
rect 194952 209585 197002 210287
rect 194952 208373 197002 209095
rect 194952 207161 197002 207883
rect 194952 205949 197002 206671
rect 194952 204737 197002 205459
rect 194952 203525 197002 204247
rect 194952 202313 197002 203035
rect 194952 201101 197002 201823
rect 194952 199889 197002 200611
rect 194952 198677 197002 199399
rect 194952 197465 197002 198187
rect 194952 196253 197002 196975
rect 194952 195041 197002 195763
rect 194952 193829 197002 194551
rect 194952 192617 197002 193339
rect 194952 191405 197002 192127
rect 194952 190193 197002 190915
rect 194952 188981 197002 189703
rect 194952 187769 197002 188491
rect 194952 186557 197002 187279
rect 194952 185345 197002 186067
rect 194952 184133 197002 184855
rect 194952 182921 197002 183643
rect 194952 181709 197002 182431
rect 194952 180497 197002 181219
rect 194952 179285 197002 180007
rect 194952 178073 197002 178795
rect 194952 176861 197002 177583
rect 194952 175649 197002 176371
rect 194952 174437 197002 175159
rect 194952 173225 197002 173947
rect 194952 172013 197002 172735
rect 194952 170630 197002 171523
rect 194952 166524 197002 170027
rect 194952 162330 197002 165136
rect 194952 159200 197002 161629
rect 194952 155404 197002 157348
rect 194952 152851 197002 154481
rect 194952 150397 197002 151720
rect 194952 105228 197002 149508
rect 194952 102748 197002 103328
rect 194952 100378 197002 100698
rect 194952 97672 197002 98328
rect 194952 95302 197002 95622
rect 194952 92672 197002 93252
rect 194952 75400 197002 90772
rect 197322 387228 199372 390292
rect 197322 384748 199372 385328
rect 197322 382378 199372 382698
rect 197322 379672 199372 380328
rect 197322 377302 199372 377622
rect 197322 374672 199372 375252
rect 197322 249581 199372 372772
rect 197322 248369 199372 249071
rect 197322 247157 199372 247859
rect 197322 245945 199372 246647
rect 197322 244733 199372 245435
rect 197322 243521 199372 244223
rect 197322 242309 199372 243011
rect 197322 241097 199372 241799
rect 197322 239885 199372 240587
rect 197322 238673 199372 239375
rect 197322 237461 199372 238163
rect 197322 236249 199372 236951
rect 197322 235037 199372 235739
rect 197322 233825 199372 234527
rect 197322 232613 199372 233315
rect 197322 231401 199372 232103
rect 197322 230189 199372 230891
rect 197322 228977 199372 229679
rect 197322 227765 199372 228467
rect 197322 226553 199372 227255
rect 197322 225341 199372 226043
rect 197322 224129 199372 224831
rect 197322 222917 199372 223619
rect 197322 221705 199372 222407
rect 197322 220493 199372 221195
rect 197322 219281 199372 219983
rect 197322 218069 199372 218771
rect 197322 216857 199372 217559
rect 197322 215645 199372 216347
rect 197322 214433 199372 215135
rect 197322 213221 199372 213923
rect 197322 212009 199372 212711
rect 197322 210797 199372 211499
rect 197322 209585 199372 210287
rect 197322 208373 199372 209095
rect 197322 207161 199372 207883
rect 197322 205949 199372 206671
rect 197322 204737 199372 205459
rect 197322 203525 199372 204247
rect 197322 202313 199372 203035
rect 197322 201101 199372 201823
rect 197322 199889 199372 200611
rect 197322 198677 199372 199399
rect 197322 197465 199372 198187
rect 197322 196253 199372 196975
rect 197322 195041 199372 195763
rect 197322 193829 199372 194551
rect 197322 192617 199372 193339
rect 197322 191405 199372 192127
rect 197322 190193 199372 190915
rect 197322 188981 199372 189703
rect 197322 187769 199372 188491
rect 197322 186557 199372 187279
rect 197322 185345 199372 186067
rect 197322 184133 199372 184855
rect 197322 182921 199372 183643
rect 197322 181709 199372 182431
rect 197322 180497 199372 181219
rect 197322 179285 199372 180007
rect 197322 178073 199372 178795
rect 197322 176861 199372 177583
rect 197322 175649 199372 176371
rect 197322 174437 199372 175159
rect 197322 173225 199372 173947
rect 197322 172013 199372 172735
rect 197322 170630 199372 171523
rect 197322 166524 199372 170027
rect 197322 162330 199372 165136
rect 197322 159200 199372 161629
rect 197322 155404 199372 157348
rect 197322 152851 199372 154481
rect 197322 150397 199372 151720
rect 197322 105228 199372 149508
rect 197322 102748 199372 103328
rect 197322 100378 199372 100698
rect 197322 97672 199372 98328
rect 197322 95302 199372 95622
rect 197322 92672 199372 93252
rect 197322 75400 199372 90772
rect 200028 387228 202078 390292
rect 200028 384748 202078 385328
rect 200028 382378 202078 382698
rect 200028 379672 202078 380328
rect 200028 377302 202078 377622
rect 200028 374672 202078 375252
rect 200028 249581 202078 372772
rect 200028 248369 202078 249071
rect 200028 247157 202078 247859
rect 200028 245945 202078 246647
rect 200028 244733 202078 245435
rect 200028 243521 202078 244223
rect 200028 242309 202078 243011
rect 200028 241097 202078 241799
rect 200028 239885 202078 240587
rect 200028 238673 202078 239375
rect 200028 237461 202078 238163
rect 200028 236249 202078 236951
rect 200028 235037 202078 235739
rect 200028 233825 202078 234527
rect 200028 232613 202078 233315
rect 200028 231401 202078 232103
rect 200028 230189 202078 230891
rect 200028 228977 202078 229679
rect 200028 227765 202078 228467
rect 200028 226553 202078 227255
rect 200028 225341 202078 226043
rect 200028 224129 202078 224831
rect 200028 222917 202078 223619
rect 200028 221705 202078 222407
rect 200028 220493 202078 221195
rect 200028 219281 202078 219983
rect 200028 218069 202078 218771
rect 200028 216857 202078 217559
rect 200028 215645 202078 216347
rect 200028 214433 202078 215135
rect 200028 213221 202078 213923
rect 200028 212009 202078 212711
rect 200028 210797 202078 211499
rect 200028 209585 202078 210287
rect 200028 208373 202078 209095
rect 200028 207161 202078 207883
rect 200028 205949 202078 206671
rect 200028 204737 202078 205459
rect 200028 203525 202078 204247
rect 200028 202313 202078 203035
rect 200028 201101 202078 201823
rect 200028 199889 202078 200611
rect 200028 198677 202078 199399
rect 200028 197465 202078 198187
rect 200028 196253 202078 196975
rect 200028 195041 202078 195763
rect 200028 193829 202078 194551
rect 200028 192617 202078 193339
rect 200028 191405 202078 192127
rect 200028 190193 202078 190915
rect 200028 188981 202078 189703
rect 200028 187769 202078 188491
rect 200028 186557 202078 187279
rect 200028 185345 202078 186067
rect 200028 184133 202078 184855
rect 200028 182921 202078 183643
rect 200028 181709 202078 182431
rect 200028 180497 202078 181219
rect 200028 179285 202078 180007
rect 200028 178073 202078 178795
rect 200028 176861 202078 177583
rect 200028 175649 202078 176371
rect 200028 174437 202078 175159
rect 200028 173225 202078 173947
rect 200028 172013 202078 172735
rect 200028 170630 202078 171523
rect 200028 166524 202078 170027
rect 200028 162330 202078 165136
rect 200028 159200 202078 161629
rect 200028 155404 202078 157348
rect 200028 152851 202078 154481
rect 200028 150397 202078 151720
rect 200028 105228 202078 149508
rect 200028 102748 202078 103328
rect 200028 100378 202078 100698
rect 200028 97672 202078 98328
rect 200028 95302 202078 95622
rect 200028 92672 202078 93252
rect 200028 75400 202078 90772
rect 202398 387228 204448 390292
rect 202398 384748 204448 385328
rect 202398 382378 204448 382698
rect 202398 379672 204448 380328
rect 202398 377302 204448 377622
rect 202398 374672 204448 375252
rect 202398 249581 204448 372772
rect 202398 248369 204448 249071
rect 202398 247157 204448 247859
rect 202398 245945 204448 246647
rect 202398 244733 204448 245435
rect 202398 243521 204448 244223
rect 202398 242309 204448 243011
rect 202398 241097 204448 241799
rect 202398 239885 204448 240587
rect 202398 238673 204448 239375
rect 202398 237461 204448 238163
rect 202398 236249 204448 236951
rect 202398 235037 204448 235739
rect 202398 233825 204448 234527
rect 202398 232613 204448 233315
rect 202398 231401 204448 232103
rect 202398 230189 204448 230891
rect 202398 228977 204448 229679
rect 202398 227765 204448 228467
rect 202398 226553 204448 227255
rect 202398 225341 204448 226043
rect 202398 224129 204448 224831
rect 202398 222917 204448 223619
rect 202398 221705 204448 222407
rect 202398 220493 204448 221195
rect 202398 219281 204448 219983
rect 202398 218069 204448 218771
rect 202398 216857 204448 217559
rect 202398 215645 204448 216347
rect 202398 214433 204448 215135
rect 202398 213221 204448 213923
rect 202398 212009 204448 212711
rect 202398 210797 204448 211499
rect 202398 209585 204448 210287
rect 202398 208373 204448 209095
rect 202398 207161 204448 207883
rect 202398 205949 204448 206671
rect 202398 204737 204448 205459
rect 202398 203525 204448 204247
rect 202398 202313 204448 203035
rect 202398 201101 204448 201823
rect 202398 199889 204448 200611
rect 202398 198677 204448 199399
rect 202398 197465 204448 198187
rect 202398 196253 204448 196975
rect 202398 195041 204448 195763
rect 202398 193829 204448 194551
rect 202398 192617 204448 193339
rect 202398 191405 204448 192127
rect 202398 190193 204448 190915
rect 202398 188981 204448 189703
rect 202398 187769 204448 188491
rect 202398 186557 204448 187279
rect 202398 185345 204448 186067
rect 202398 184133 204448 184855
rect 202398 182921 204448 183643
rect 202398 181709 204448 182431
rect 202398 180497 204448 181219
rect 202398 179285 204448 180007
rect 202398 178073 204448 178795
rect 202398 176861 204448 177583
rect 202398 175649 204448 176371
rect 202398 174437 204448 175159
rect 202398 173225 204448 173947
rect 202398 172013 204448 172735
rect 202398 170630 204448 171523
rect 202398 166524 204448 170027
rect 202398 162330 204448 165136
rect 202398 159200 204448 161629
rect 202398 155404 204448 157348
rect 202398 152851 204448 154481
rect 202398 150397 204448 151720
rect 202398 105228 204448 149508
rect 202398 102748 204448 103328
rect 202398 100378 204448 100698
rect 202398 97672 204448 98328
rect 202398 95302 204448 95622
rect 202398 92672 204448 93252
rect 202398 75400 204448 90772
rect 205028 387228 206851 390292
rect 205028 384748 206851 385328
rect 205028 382378 206851 382698
rect 205028 379672 206851 380328
rect 205028 377302 206851 377622
rect 205028 374672 206851 375252
rect 205028 249581 206851 372772
rect 205028 248369 206851 249071
rect 205028 247157 206851 247859
rect 205028 245945 206851 246647
rect 205028 244733 206851 245435
rect 205028 243521 206851 244223
rect 205028 242309 206851 243011
rect 205028 241097 206851 241799
rect 205028 239885 206851 240587
rect 205028 238673 206851 239375
rect 205028 237461 206851 238163
rect 205028 236249 206851 236951
rect 205028 235037 206851 235739
rect 205028 233825 206851 234527
rect 205028 232613 206851 233315
rect 205028 231401 206851 232103
rect 205028 230189 206851 230891
rect 205028 228977 206851 229679
rect 205028 227765 206851 228467
rect 205028 226553 206851 227255
rect 205028 225341 206851 226043
rect 205028 224129 206851 224831
rect 205028 222917 206851 223619
rect 205028 221705 206851 222407
rect 205028 220493 206851 221195
rect 205028 219281 206851 219983
rect 205028 218069 206851 218771
rect 205028 216857 206851 217559
rect 205028 215645 206851 216347
rect 205028 214433 206851 215135
rect 205028 213221 206851 213923
rect 205028 212009 206851 212711
rect 205028 210797 206851 211499
rect 205028 209585 206851 210287
rect 205028 208373 206851 209095
rect 205028 207161 206851 207883
rect 205028 205949 206851 206671
rect 205028 204737 206851 205459
rect 205028 203525 206851 204247
rect 205028 202313 206851 203035
rect 205028 201101 206851 201823
rect 205028 199889 206851 200611
rect 205028 198677 206851 199399
rect 205028 197465 206851 198187
rect 205028 196253 206851 196975
rect 205028 195041 206851 195763
rect 205028 193829 206851 194551
rect 205028 192617 206851 193339
rect 205028 191405 206851 192127
rect 205028 190193 206851 190915
rect 205028 188981 206851 189703
rect 205028 187769 206851 188491
rect 205028 186557 206851 187279
rect 205028 185345 206851 186067
rect 205028 184133 206851 184855
rect 205028 182921 206851 183643
rect 205028 181709 206851 182431
rect 205028 180497 206851 181219
rect 205028 179285 206851 180007
rect 205028 178073 206851 178795
rect 205028 176861 206851 177583
rect 205028 175649 206851 176371
rect 205028 174437 206851 175159
rect 205028 173225 206851 173947
rect 205028 172013 206851 172735
rect 205028 170630 206851 171523
rect 205028 166524 206851 170027
rect 205028 162330 206851 165136
rect 205028 159200 206851 161629
rect 205028 155404 206851 157348
rect 205028 152851 206851 154481
rect 205028 150397 206851 151720
rect 205028 105228 206851 149508
rect 205028 102748 206851 103328
rect 205028 100378 206851 100698
rect 205028 97672 206851 98328
rect 205028 95302 206851 95622
rect 205028 92672 206851 93252
rect 205028 75400 206851 90772
rect 218272 250360 220172 400972
rect 218272 248971 220172 249660
rect 218272 247759 220172 248481
rect 218272 246547 220172 247269
rect 218272 245335 220172 246057
rect 218272 244123 220172 244845
rect 218272 242911 220172 243633
rect 218272 241699 220172 242421
rect 218272 240487 220172 241209
rect 218272 239275 220172 239997
rect 218272 238063 220172 238785
rect 218272 236851 220172 237573
rect 218272 235639 220172 236361
rect 218272 234427 220172 235149
rect 218272 233215 220172 233937
rect 218272 232003 220172 232725
rect 218272 230791 220172 231513
rect 218272 229579 220172 230301
rect 218272 228367 220172 229089
rect 218272 227155 220172 227877
rect 218272 225943 220172 226665
rect 218272 224731 220172 225453
rect 218272 223519 220172 224241
rect 218272 222307 220172 223029
rect 218272 221095 220172 221817
rect 218272 219883 220172 220605
rect 218272 218671 220172 219393
rect 218272 217459 220172 218181
rect 218272 216247 220172 216969
rect 218272 215035 220172 215757
rect 218272 213823 220172 214545
rect 218272 212611 220172 213333
rect 218272 211576 220172 212121
rect 218272 210187 220172 210876
rect 218272 208975 220172 209697
rect 218272 207763 220172 208485
rect 218272 206551 220172 207273
rect 218272 205339 220172 206061
rect 218272 204127 220172 204849
rect 218272 202915 220172 203637
rect 218272 201703 220172 202425
rect 218272 200491 220172 201213
rect 218272 199279 220172 200001
rect 218272 198067 220172 198789
rect 218272 196855 220172 197577
rect 218272 195643 220172 196365
rect 218272 194431 220172 195153
rect 218272 193219 220172 193941
rect 218272 192007 220172 192729
rect 218272 190795 220172 191517
rect 218272 189583 220172 190305
rect 218272 188371 220172 189093
rect 218272 187159 220172 187881
rect 218272 185947 220172 186669
rect 218272 184735 220172 185457
rect 218272 183523 220172 184245
rect 218272 182311 220172 183033
rect 218272 181099 220172 181821
rect 218272 179887 220172 180609
rect 218272 178675 220172 179397
rect 218272 177463 220172 178185
rect 218272 176251 220172 176973
rect 218272 175039 220172 175761
rect 218272 173827 220172 174549
rect 218272 172615 220172 173337
rect 218272 171403 220172 172125
rect 218272 169740 220172 170913
rect 218272 163429 220172 166792
rect 218272 161308 220172 162728
rect 218272 157222 220172 159399
rect 218272 154018 220172 155760
rect 218272 151628 220172 153063
rect 218272 149320 220172 150599
rect 218272 133428 220172 148620
rect 218272 130948 220172 131528
rect 218272 128578 220172 128898
rect 218272 125872 220172 126528
rect 218272 123502 220172 123822
rect 218272 120872 220172 121452
rect 218272 87078 220172 118972
rect 218272 75400 220172 86550
rect 220752 415428 222802 417503
rect 220752 412948 222802 413528
rect 220752 410578 222802 410898
rect 220752 407872 222802 408528
rect 220752 405502 222802 405822
rect 220752 402872 222802 403452
rect 220752 250360 222802 400972
rect 220752 248971 222802 249660
rect 220752 247759 222802 248481
rect 220752 246547 222802 247269
rect 220752 245335 222802 246057
rect 220752 244123 222802 244845
rect 220752 242911 222802 243633
rect 220752 241699 222802 242421
rect 220752 240487 222802 241209
rect 220752 239275 222802 239997
rect 220752 238063 222802 238785
rect 220752 236851 222802 237573
rect 220752 235639 222802 236361
rect 220752 234427 222802 235149
rect 220752 233215 222802 233937
rect 220752 232003 222802 232725
rect 220752 230791 222802 231513
rect 220752 229579 222802 230301
rect 220752 228367 222802 229089
rect 220752 227155 222802 227877
rect 220752 225943 222802 226665
rect 220752 224731 222802 225453
rect 220752 223519 222802 224241
rect 220752 222307 222802 223029
rect 220752 221095 222802 221817
rect 220752 219883 222802 220605
rect 220752 218671 222802 219393
rect 220752 217459 222802 218181
rect 220752 216247 222802 216969
rect 220752 215035 222802 215757
rect 220752 213823 222802 214545
rect 220752 212611 222802 213333
rect 220752 211576 222802 212121
rect 220752 210187 222802 210876
rect 220752 208975 222802 209697
rect 220752 207763 222802 208485
rect 220752 206551 222802 207273
rect 220752 205339 222802 206061
rect 220752 204127 222802 204849
rect 220752 202915 222802 203637
rect 220752 201703 222802 202425
rect 220752 200491 222802 201213
rect 220752 199279 222802 200001
rect 220752 198067 222802 198789
rect 220752 196855 222802 197577
rect 220752 195643 222802 196365
rect 220752 194431 222802 195153
rect 220752 193219 222802 193941
rect 220752 192007 222802 192729
rect 220752 190795 222802 191517
rect 220752 189583 222802 190305
rect 220752 188371 222802 189093
rect 220752 187159 222802 187881
rect 220752 185947 222802 186669
rect 220752 184735 222802 185457
rect 220752 183523 222802 184245
rect 220752 182311 222802 183033
rect 220752 181099 222802 181821
rect 220752 179887 222802 180609
rect 220752 178675 222802 179397
rect 220752 177463 222802 178185
rect 220752 176251 222802 176973
rect 220752 175039 222802 175761
rect 220752 173827 222802 174549
rect 220752 172615 222802 173337
rect 220752 171403 222802 172125
rect 220752 169740 222802 170913
rect 220752 163429 222802 166792
rect 220752 161308 222802 162728
rect 220752 157222 222802 159399
rect 220752 154018 222802 155760
rect 220752 151628 222802 153063
rect 220752 149320 222802 150599
rect 220752 133428 222802 148620
rect 220752 130948 222802 131528
rect 220752 128578 222802 128898
rect 220752 125872 222802 126528
rect 220752 123502 222802 123822
rect 220752 120872 222802 121452
rect 220752 75400 222802 118972
rect 223122 415428 225172 417503
rect 223122 412948 225172 413528
rect 223122 410578 225172 410898
rect 223122 407872 225172 408528
rect 223122 405502 225172 405822
rect 223122 402872 225172 403452
rect 223122 250360 225172 400972
rect 223122 248971 225172 249660
rect 223122 247759 225172 248481
rect 223122 246547 225172 247269
rect 223122 245335 225172 246057
rect 223122 244123 225172 244845
rect 223122 242911 225172 243633
rect 223122 241699 225172 242421
rect 223122 240487 225172 241209
rect 223122 239275 225172 239997
rect 223122 238063 225172 238785
rect 223122 236851 225172 237573
rect 223122 235639 225172 236361
rect 223122 234427 225172 235149
rect 223122 233215 225172 233937
rect 223122 232003 225172 232725
rect 223122 230791 225172 231513
rect 223122 229579 225172 230301
rect 223122 228367 225172 229089
rect 223122 227155 225172 227877
rect 223122 225943 225172 226665
rect 223122 224731 225172 225453
rect 223122 223519 225172 224241
rect 223122 222307 225172 223029
rect 223122 221095 225172 221817
rect 223122 219883 225172 220605
rect 223122 218671 225172 219393
rect 223122 217459 225172 218181
rect 223122 216247 225172 216969
rect 223122 215035 225172 215757
rect 223122 213823 225172 214545
rect 223122 212611 225172 213333
rect 223122 211576 225172 212121
rect 223122 210187 225172 210876
rect 223122 208975 225172 209697
rect 223122 207763 225172 208485
rect 223122 206551 225172 207273
rect 223122 205339 225172 206061
rect 223122 204127 225172 204849
rect 223122 202915 225172 203637
rect 223122 201703 225172 202425
rect 223122 200491 225172 201213
rect 223122 199279 225172 200001
rect 223122 198067 225172 198789
rect 223122 196855 225172 197577
rect 223122 195643 225172 196365
rect 223122 194431 225172 195153
rect 223122 193219 225172 193941
rect 223122 192007 225172 192729
rect 223122 190795 225172 191517
rect 223122 189583 225172 190305
rect 223122 188371 225172 189093
rect 223122 187159 225172 187881
rect 223122 185947 225172 186669
rect 223122 184735 225172 185457
rect 223122 183523 225172 184245
rect 223122 182311 225172 183033
rect 223122 181099 225172 181821
rect 223122 179887 225172 180609
rect 223122 178675 225172 179397
rect 223122 177463 225172 178185
rect 223122 176251 225172 176973
rect 223122 175039 225172 175761
rect 223122 173827 225172 174549
rect 223122 172615 225172 173337
rect 223122 171403 225172 172125
rect 223122 169740 225172 170913
rect 223122 163429 225172 166792
rect 223122 161308 225172 162728
rect 223122 157222 225172 159399
rect 223122 154018 225172 155760
rect 223122 151628 225172 153063
rect 223122 149320 225172 150599
rect 223122 133428 225172 148620
rect 223122 130948 225172 131528
rect 223122 128578 225172 128898
rect 223122 125872 225172 126528
rect 223122 123502 225172 123822
rect 223122 120872 225172 121452
rect 223122 75400 225172 118972
rect 225828 415428 227878 417503
rect 225828 412948 227878 413528
rect 225828 410578 227878 410898
rect 225828 407872 227878 408528
rect 225828 405502 227878 405822
rect 225828 402872 227878 403452
rect 225828 250360 227878 400972
rect 225828 248971 227878 249660
rect 225828 247759 227878 248481
rect 225828 246547 227878 247269
rect 225828 245335 227878 246057
rect 225828 244123 227878 244845
rect 225828 242911 227878 243633
rect 225828 241699 227878 242421
rect 225828 240487 227878 241209
rect 225828 239275 227878 239997
rect 225828 238063 227878 238785
rect 225828 236851 227878 237573
rect 225828 235639 227878 236361
rect 225828 234427 227878 235149
rect 225828 233215 227878 233937
rect 225828 232003 227878 232725
rect 225828 230791 227878 231513
rect 225828 229579 227878 230301
rect 225828 228367 227878 229089
rect 225828 227155 227878 227877
rect 225828 225943 227878 226665
rect 225828 224731 227878 225453
rect 225828 223519 227878 224241
rect 225828 222307 227878 223029
rect 225828 221095 227878 221817
rect 225828 219883 227878 220605
rect 225828 218671 227878 219393
rect 225828 217459 227878 218181
rect 225828 216247 227878 216969
rect 225828 215035 227878 215757
rect 225828 213823 227878 214545
rect 225828 212611 227878 213333
rect 225828 211576 227878 212121
rect 225828 210187 227878 210876
rect 225828 208975 227878 209697
rect 225828 207763 227878 208485
rect 225828 206551 227878 207273
rect 225828 205339 227878 206061
rect 225828 204127 227878 204849
rect 225828 202915 227878 203637
rect 225828 201703 227878 202425
rect 225828 200491 227878 201213
rect 225828 199279 227878 200001
rect 225828 198067 227878 198789
rect 225828 196855 227878 197577
rect 225828 195643 227878 196365
rect 225828 194431 227878 195153
rect 225828 193219 227878 193941
rect 225828 192007 227878 192729
rect 225828 190795 227878 191517
rect 225828 189583 227878 190305
rect 225828 188371 227878 189093
rect 225828 187159 227878 187881
rect 225828 185947 227878 186669
rect 225828 184735 227878 185457
rect 225828 183523 227878 184245
rect 225828 182311 227878 183033
rect 225828 181099 227878 181821
rect 225828 179887 227878 180609
rect 225828 178675 227878 179397
rect 225828 177463 227878 178185
rect 225828 176251 227878 176973
rect 225828 175039 227878 175761
rect 225828 173827 227878 174549
rect 225828 172615 227878 173337
rect 225828 171403 227878 172125
rect 225828 169740 227878 170913
rect 225828 163429 227878 166792
rect 225828 161308 227878 162728
rect 225828 157222 227878 159399
rect 225828 154018 227878 155760
rect 225828 151628 227878 153063
rect 225828 149320 227878 150599
rect 225828 133428 227878 148620
rect 225828 130948 227878 131528
rect 225828 128578 227878 128898
rect 225828 125872 227878 126528
rect 225828 123502 227878 123822
rect 225828 120872 227878 121452
rect 225828 75400 227878 118972
rect 228198 415428 230248 417503
rect 228198 412948 230248 413528
rect 228198 410578 230248 410898
rect 228198 407872 230248 408528
rect 228198 405502 230248 405822
rect 228198 402872 230248 403452
rect 228198 250360 230248 400972
rect 228198 248971 230248 249660
rect 228198 247759 230248 248481
rect 228198 246547 230248 247269
rect 228198 245335 230248 246057
rect 228198 244123 230248 244845
rect 228198 242911 230248 243633
rect 228198 241699 230248 242421
rect 228198 240487 230248 241209
rect 228198 239275 230248 239997
rect 228198 238063 230248 238785
rect 228198 236851 230248 237573
rect 228198 235639 230248 236361
rect 228198 234427 230248 235149
rect 228198 233215 230248 233937
rect 228198 232003 230248 232725
rect 228198 230791 230248 231513
rect 228198 229579 230248 230301
rect 228198 228367 230248 229089
rect 228198 227155 230248 227877
rect 228198 225943 230248 226665
rect 228198 224731 230248 225453
rect 228198 223519 230248 224241
rect 228198 222307 230248 223029
rect 228198 221095 230248 221817
rect 228198 219883 230248 220605
rect 228198 218671 230248 219393
rect 228198 217459 230248 218181
rect 228198 216247 230248 216969
rect 228198 215035 230248 215757
rect 228198 213823 230248 214545
rect 228198 212611 230248 213333
rect 228198 211576 230248 212121
rect 228198 210187 230248 210876
rect 228198 208975 230248 209697
rect 228198 207763 230248 208485
rect 228198 206551 230248 207273
rect 228198 205339 230248 206061
rect 228198 204127 230248 204849
rect 228198 202915 230248 203637
rect 228198 201703 230248 202425
rect 228198 200491 230248 201213
rect 228198 199279 230248 200001
rect 228198 198067 230248 198789
rect 228198 196855 230248 197577
rect 228198 195643 230248 196365
rect 228198 194431 230248 195153
rect 228198 193219 230248 193941
rect 228198 192007 230248 192729
rect 228198 190795 230248 191517
rect 228198 189583 230248 190305
rect 228198 188371 230248 189093
rect 228198 187159 230248 187881
rect 228198 185947 230248 186669
rect 228198 184735 230248 185457
rect 228198 183523 230248 184245
rect 228198 182311 230248 183033
rect 228198 181099 230248 181821
rect 228198 179887 230248 180609
rect 228198 178675 230248 179397
rect 228198 177463 230248 178185
rect 228198 176251 230248 176973
rect 228198 175039 230248 175761
rect 228198 173827 230248 174549
rect 228198 172615 230248 173337
rect 228198 171403 230248 172125
rect 228198 169740 230248 170913
rect 228198 163429 230248 166792
rect 228198 161308 230248 162728
rect 228198 157222 230248 159399
rect 228198 154018 230248 155760
rect 228198 151628 230248 153063
rect 228198 149320 230248 150599
rect 228198 133428 230248 148620
rect 228198 130948 230248 131528
rect 228198 128578 230248 128898
rect 228198 125872 230248 126528
rect 228198 123502 230248 123822
rect 228198 120872 230248 121452
rect 228198 75400 230248 118972
rect 230828 415428 232655 417503
rect 230828 412948 232655 413528
rect 230828 410578 232655 410898
rect 230828 407872 232655 408528
rect 230828 405502 232655 405822
rect 230828 402872 232655 403452
rect 230828 250360 232655 400972
rect 230828 248971 232655 249660
rect 230828 247759 232655 248481
rect 230828 246547 232655 247269
rect 230828 245335 232655 246057
rect 230828 244123 232655 244845
rect 230828 242911 232655 243633
rect 230828 241699 232655 242421
rect 230828 240487 232655 241209
rect 230828 239275 232655 239997
rect 230828 238063 232655 238785
rect 230828 236851 232655 237573
rect 230828 235639 232655 236361
rect 230828 234427 232655 235149
rect 230828 233215 232655 233937
rect 230828 232003 232655 232725
rect 230828 230791 232655 231513
rect 230828 229579 232655 230301
rect 230828 228367 232655 229089
rect 230828 227155 232655 227877
rect 230828 225943 232655 226665
rect 230828 224731 232655 225453
rect 230828 223519 232655 224241
rect 230828 222307 232655 223029
rect 230828 221095 232655 221817
rect 230828 219883 232655 220605
rect 230828 218671 232655 219393
rect 230828 217459 232655 218181
rect 230828 216247 232655 216969
rect 230828 215035 232655 215757
rect 230828 213823 232655 214545
rect 230828 212611 232655 213333
rect 230828 211576 232655 212121
rect 230828 210187 232655 210876
rect 230828 208975 232655 209697
rect 230828 207763 232655 208485
rect 230828 206551 232655 207273
rect 230828 205339 232655 206061
rect 230828 204127 232655 204849
rect 230828 202915 232655 203637
rect 230828 201703 232655 202425
rect 230828 200491 232655 201213
rect 230828 199279 232655 200001
rect 230828 198067 232655 198789
rect 230828 196855 232655 197577
rect 230828 195643 232655 196365
rect 230828 194431 232655 195153
rect 230828 193219 232655 193941
rect 230828 192007 232655 192729
rect 230828 190795 232655 191517
rect 230828 189583 232655 190305
rect 230828 188371 232655 189093
rect 230828 187159 232655 187881
rect 230828 185947 232655 186669
rect 230828 184735 232655 185457
rect 230828 183523 232655 184245
rect 230828 182311 232655 183033
rect 230828 181099 232655 181821
rect 230828 179887 232655 180609
rect 230828 178675 232655 179397
rect 230828 177463 232655 178185
rect 230828 176251 232655 176973
rect 230828 175039 232655 175761
rect 230828 173827 232655 174549
rect 230828 172615 232655 173337
rect 230828 171403 232655 172125
rect 230828 169740 232655 170913
rect 230828 163429 232655 166792
rect 230828 161308 232655 162728
rect 230828 157222 232655 159399
rect 230828 154018 232655 155760
rect 230828 151628 232655 153063
rect 553672 387228 555572 430800
rect 553672 384748 555572 385328
rect 553672 382378 555572 382698
rect 553672 379672 555572 380328
rect 553672 377302 555572 377622
rect 553672 374672 555572 375252
rect 553672 190904 555572 372772
rect 553672 189692 555572 190394
rect 553672 188480 555572 189202
rect 553672 187268 555572 187990
rect 553672 186056 555572 186778
rect 553672 184844 555572 185566
rect 553672 183632 555572 184354
rect 553672 182420 555572 183142
rect 553672 181208 555572 181930
rect 553672 179996 555572 180718
rect 553672 178784 555572 179506
rect 553672 177572 555572 178294
rect 553672 176360 555572 177082
rect 553672 175148 555572 175870
rect 553672 173936 555572 174658
rect 553672 172724 555572 173446
rect 553672 171512 555572 172234
rect 553672 170129 555572 171022
rect 553672 166023 555572 169526
rect 553672 161829 555572 164635
rect 553672 158699 555572 161128
rect 553672 154903 555572 156847
rect 553672 152350 555572 153980
rect 230828 149320 232655 150599
rect 230828 133428 232655 148620
rect 230828 130948 232655 131528
rect 230828 128578 232655 128898
rect 230828 125872 232655 126528
rect 230828 123502 232655 123822
rect 230828 120872 232655 121452
rect 230828 75400 232655 118972
rect 327021 149232 327835 150683
rect 327021 105228 327835 149098
rect 327021 102748 327835 103328
rect 327021 100378 327835 100698
rect 327021 97672 327835 98328
rect 327021 95302 327835 95622
rect 327021 92672 327835 93252
rect 327021 90489 327835 90772
rect 328649 150030 329463 150683
rect 328649 133428 329463 149896
rect 328649 130948 329463 131528
rect 328649 128578 329463 128898
rect 328649 125872 329463 126528
rect 328649 123502 329463 123822
rect 328649 120872 329463 121452
rect 328649 90489 329463 118972
rect 459446 150332 460246 150444
rect 459446 133428 460246 150035
rect 459446 130948 460246 131528
rect 459446 128578 460246 128898
rect 459446 125872 460246 126528
rect 459446 123502 460246 123822
rect 459446 120872 460246 121452
rect 459446 90126 460246 118972
rect 460979 149711 461779 150405
rect 460979 105228 461779 149414
rect 460979 102748 461779 103328
rect 460979 100378 461779 100698
rect 460979 97672 461779 98328
rect 460979 95302 461779 95622
rect 460979 92672 461779 93252
rect 460979 90169 461779 90772
rect 553672 149896 555572 151219
rect 553672 105228 555572 149007
rect 553672 102748 555572 103328
rect 553672 100378 555572 100698
rect 553672 97672 555572 98328
rect 553672 95302 555572 95622
rect 553672 92672 555572 93252
rect 553672 89056 555572 90772
rect 556152 387228 558202 430800
rect 556152 384748 558202 385328
rect 556152 382378 558202 382698
rect 556152 379672 558202 380328
rect 556152 377302 558202 377622
rect 556152 374672 558202 375252
rect 556152 190904 558202 372772
rect 556152 189692 558202 190394
rect 556152 188480 558202 189202
rect 556152 187268 558202 187990
rect 556152 186056 558202 186778
rect 556152 184844 558202 185566
rect 556152 183632 558202 184354
rect 556152 182420 558202 183142
rect 556152 181208 558202 181930
rect 556152 179996 558202 180718
rect 556152 178784 558202 179506
rect 556152 177572 558202 178294
rect 556152 176360 558202 177082
rect 556152 175148 558202 175870
rect 556152 173936 558202 174658
rect 556152 172724 558202 173446
rect 556152 171512 558202 172234
rect 556152 170129 558202 171022
rect 556152 166023 558202 169526
rect 556152 161829 558202 164635
rect 556152 158699 558202 161128
rect 556152 154903 558202 156847
rect 556152 152350 558202 153980
rect 556152 149896 558202 151219
rect 556152 105228 558202 149007
rect 556152 102748 558202 103328
rect 556152 100378 558202 100698
rect 556152 97672 558202 98328
rect 556152 95302 558202 95622
rect 556152 92672 558202 93252
rect 556152 89056 558202 90772
rect 558522 387228 560572 430800
rect 558522 384748 560572 385328
rect 558522 382378 560572 382698
rect 558522 379672 560572 380328
rect 558522 377302 560572 377622
rect 558522 374672 560572 375252
rect 558522 190904 560572 372772
rect 558522 189692 560572 190394
rect 558522 188480 560572 189202
rect 558522 187268 560572 187990
rect 558522 186056 560572 186778
rect 558522 184844 560572 185566
rect 558522 183632 560572 184354
rect 558522 182420 560572 183142
rect 558522 181208 560572 181930
rect 558522 179996 560572 180718
rect 558522 178784 560572 179506
rect 558522 177572 560572 178294
rect 558522 176360 560572 177082
rect 558522 175148 560572 175870
rect 558522 173936 560572 174658
rect 558522 172724 560572 173446
rect 558522 171512 560572 172234
rect 558522 170129 560572 171022
rect 558522 166023 560572 169526
rect 558522 161829 560572 164635
rect 558522 158699 560572 161128
rect 558522 154903 560572 156847
rect 558522 152350 560572 153980
rect 558522 149896 560572 151219
rect 558522 105228 560572 149007
rect 558522 102748 560572 103328
rect 558522 100378 560572 100698
rect 558522 97672 560572 98328
rect 558522 95302 560572 95622
rect 558522 92672 560572 93252
rect 558522 89056 560572 90772
rect 561228 387228 563278 430800
rect 561228 384748 563278 385328
rect 561228 382378 563278 382698
rect 561228 379672 563278 380328
rect 561228 377302 563278 377622
rect 561228 374672 563278 375252
rect 561228 190904 563278 372772
rect 561228 189692 563278 190394
rect 561228 188480 563278 189202
rect 561228 187268 563278 187990
rect 561228 186056 563278 186778
rect 561228 184844 563278 185566
rect 561228 183632 563278 184354
rect 561228 182420 563278 183142
rect 561228 181208 563278 181930
rect 561228 179996 563278 180718
rect 561228 178784 563278 179506
rect 561228 177572 563278 178294
rect 561228 176360 563278 177082
rect 561228 175148 563278 175870
rect 561228 173936 563278 174658
rect 561228 172724 563278 173446
rect 561228 171512 563278 172234
rect 561228 170129 563278 171022
rect 561228 166023 563278 169526
rect 561228 161829 563278 164635
rect 561228 158699 563278 161128
rect 561228 154903 563278 156847
rect 561228 152350 563278 153980
rect 561228 149896 563278 151219
rect 561228 105228 563278 149007
rect 561228 102748 563278 103328
rect 561228 100378 563278 100698
rect 561228 97672 563278 98328
rect 561228 95302 563278 95622
rect 561228 92672 563278 93252
rect 561228 89056 563278 90772
rect 563598 387228 565648 430800
rect 563598 384748 565648 385328
rect 563598 382378 565648 382698
rect 563598 379672 565648 380328
rect 563598 377302 565648 377622
rect 563598 374672 565648 375252
rect 563598 190904 565648 372772
rect 563598 189692 565648 190394
rect 563598 188480 565648 189202
rect 563598 187268 565648 187990
rect 563598 186056 565648 186778
rect 563598 184844 565648 185566
rect 563598 183632 565648 184354
rect 563598 182420 565648 183142
rect 563598 181208 565648 181930
rect 563598 179996 565648 180718
rect 563598 178784 565648 179506
rect 563598 177572 565648 178294
rect 563598 176360 565648 177082
rect 563598 175148 565648 175870
rect 563598 173936 565648 174658
rect 563598 172724 565648 173446
rect 563598 171512 565648 172234
rect 563598 170129 565648 171022
rect 563598 166023 565648 169526
rect 563598 161829 565648 164635
rect 563598 158699 565648 161128
rect 563598 154903 565648 156847
rect 563598 152350 565648 153980
rect 563598 149896 565648 151219
rect 563598 105228 565648 149007
rect 563598 102748 565648 103328
rect 563598 100378 565648 100698
rect 563598 97672 565648 98328
rect 563598 95302 565648 95622
rect 563598 92672 565648 93252
rect 563598 89056 565648 90772
rect 566228 387228 568128 430800
rect 566228 384748 568128 385328
rect 566228 382378 568128 382698
rect 566228 379672 568128 380328
rect 566228 377302 568128 377622
rect 566228 374672 568128 375252
rect 566228 190904 568128 372772
rect 566228 189692 568128 190394
rect 566228 188480 568128 189202
rect 566228 187268 568128 187990
rect 566228 186056 568128 186778
rect 566228 184844 568128 185566
rect 566228 183632 568128 184354
rect 566228 182420 568128 183142
rect 566228 181208 568128 181930
rect 566228 179996 568128 180718
rect 566228 178784 568128 179506
rect 566228 177572 568128 178294
rect 566228 176360 568128 177082
rect 566228 175148 568128 175870
rect 566228 173936 568128 174658
rect 566228 172724 568128 173446
rect 566228 171512 568128 172234
rect 566228 170129 568128 171022
rect 566228 166023 568128 169526
rect 566228 161829 568128 164635
rect 566228 158699 568128 161128
rect 566228 154903 568128 156847
rect 566228 152350 568128 153980
rect 566228 149896 568128 151219
rect 566228 105228 568128 149007
rect 579472 415428 581372 430800
rect 579472 412948 581372 413528
rect 579472 410578 581372 410898
rect 579472 407872 581372 408528
rect 579472 405502 581372 405822
rect 579472 402872 581372 403452
rect 579472 191683 581372 400972
rect 579472 190294 581372 190983
rect 579472 189082 581372 189804
rect 579472 187870 581372 188592
rect 579472 186658 581372 187380
rect 579472 185446 581372 186168
rect 579472 184234 581372 184956
rect 579472 183022 581372 183744
rect 579472 181810 581372 182532
rect 579472 180598 581372 181320
rect 579472 179386 581372 180108
rect 579472 178174 581372 178896
rect 579472 176962 581372 177684
rect 579472 175750 581372 176472
rect 579472 174538 581372 175260
rect 579472 173326 581372 174048
rect 579472 172114 581372 172836
rect 579472 170902 581372 171624
rect 579472 169239 581372 170412
rect 579472 162928 581372 166291
rect 579472 160807 581372 162227
rect 579472 156721 581372 158898
rect 579472 153517 581372 155259
rect 579472 151127 581372 152562
rect 579472 148819 581372 150098
rect 579472 133428 581372 148119
rect 579472 130948 581372 131528
rect 579472 128578 581372 128898
rect 579472 125872 581372 126528
rect 579472 123502 581372 123822
rect 579472 120872 581372 121452
rect 579472 116651 581372 118972
rect 581952 415428 584002 430800
rect 581952 412948 584002 413528
rect 581952 410578 584002 410898
rect 581952 407872 584002 408528
rect 581952 405502 584002 405822
rect 581952 402872 584002 403452
rect 581952 191683 584002 400972
rect 581952 190294 584002 190983
rect 581952 189082 584002 189804
rect 581952 187870 584002 188592
rect 581952 186658 584002 187380
rect 581952 185446 584002 186168
rect 581952 184234 584002 184956
rect 581952 183022 584002 183744
rect 581952 181810 584002 182532
rect 581952 180598 584002 181320
rect 581952 179386 584002 180108
rect 581952 178174 584002 178896
rect 581952 176962 584002 177684
rect 581952 175750 584002 176472
rect 581952 174538 584002 175260
rect 581952 173326 584002 174048
rect 581952 172114 584002 172836
rect 581952 170902 584002 171624
rect 581952 169239 584002 170412
rect 581952 162928 584002 166291
rect 581952 160807 584002 162227
rect 581952 156721 584002 158898
rect 581952 153517 584002 155259
rect 581952 151127 584002 152562
rect 581952 148819 584002 150098
rect 581952 133428 584002 148119
rect 581952 130948 584002 131528
rect 581952 128578 584002 128898
rect 581952 125872 584002 126528
rect 581952 123502 584002 123822
rect 581952 120872 584002 121452
rect 581952 116651 584002 118972
rect 584322 415428 586372 430800
rect 584322 412948 586372 413528
rect 584322 410578 586372 410898
rect 584322 407872 586372 408528
rect 584322 405502 586372 405822
rect 584322 402872 586372 403452
rect 584322 191683 586372 400972
rect 584322 190294 586372 190983
rect 584322 189082 586372 189804
rect 584322 187870 586372 188592
rect 584322 186658 586372 187380
rect 584322 185446 586372 186168
rect 584322 184234 586372 184956
rect 584322 183022 586372 183744
rect 584322 181810 586372 182532
rect 584322 180598 586372 181320
rect 584322 179386 586372 180108
rect 584322 178174 586372 178896
rect 584322 176962 586372 177684
rect 584322 175750 586372 176472
rect 584322 174538 586372 175260
rect 584322 173326 586372 174048
rect 584322 172114 586372 172836
rect 584322 170902 586372 171624
rect 584322 169239 586372 170412
rect 584322 162928 586372 166291
rect 584322 160807 586372 162227
rect 584322 156721 586372 158898
rect 584322 153517 586372 155259
rect 584322 151127 586372 152562
rect 584322 148819 586372 150098
rect 584322 133428 586372 148119
rect 584322 130948 586372 131528
rect 584322 128578 586372 128898
rect 584322 125872 586372 126528
rect 584322 123502 586372 123822
rect 584322 120872 586372 121452
rect 584322 116651 586372 118972
rect 587028 415428 589078 430800
rect 587028 412948 589078 413528
rect 587028 410578 589078 410898
rect 587028 407872 589078 408528
rect 587028 405502 589078 405822
rect 587028 402872 589078 403452
rect 587028 191683 589078 400972
rect 587028 190294 589078 190983
rect 587028 189082 589078 189804
rect 587028 187870 589078 188592
rect 587028 186658 589078 187380
rect 587028 185446 589078 186168
rect 587028 184234 589078 184956
rect 587028 183022 589078 183744
rect 587028 181810 589078 182532
rect 587028 180598 589078 181320
rect 587028 179386 589078 180108
rect 587028 178174 589078 178896
rect 587028 176962 589078 177684
rect 587028 175750 589078 176472
rect 587028 174538 589078 175260
rect 587028 173326 589078 174048
rect 587028 172114 589078 172836
rect 587028 170902 589078 171624
rect 587028 169239 589078 170412
rect 587028 162928 589078 166291
rect 587028 160807 589078 162227
rect 587028 156721 589078 158898
rect 587028 153517 589078 155259
rect 587028 151127 589078 152562
rect 587028 148819 589078 150098
rect 587028 133428 589078 148119
rect 587028 130948 589078 131528
rect 587028 128578 589078 128898
rect 587028 125872 589078 126528
rect 587028 123502 589078 123822
rect 587028 120872 589078 121452
rect 587028 116651 589078 118972
rect 589398 415428 591448 430800
rect 589398 412948 591448 413528
rect 589398 410578 591448 410898
rect 589398 407872 591448 408528
rect 589398 405502 591448 405822
rect 589398 402872 591448 403452
rect 589398 191683 591448 400972
rect 589398 190294 591448 190983
rect 589398 189082 591448 189804
rect 589398 187870 591448 188592
rect 589398 186658 591448 187380
rect 589398 185446 591448 186168
rect 589398 184234 591448 184956
rect 589398 183022 591448 183744
rect 589398 181810 591448 182532
rect 589398 180598 591448 181320
rect 589398 179386 591448 180108
rect 589398 178174 591448 178896
rect 589398 176962 591448 177684
rect 589398 175750 591448 176472
rect 589398 174538 591448 175260
rect 589398 173326 591448 174048
rect 589398 172114 591448 172836
rect 589398 170902 591448 171624
rect 589398 169239 591448 170412
rect 589398 162928 591448 166291
rect 589398 160807 591448 162227
rect 589398 156721 591448 158898
rect 589398 153517 591448 155259
rect 589398 151127 591448 152562
rect 589398 148819 591448 150098
rect 589398 133428 591448 148119
rect 589398 130948 591448 131528
rect 589398 128578 591448 128898
rect 589398 125872 591448 126528
rect 589398 123502 591448 123822
rect 589398 120872 591448 121452
rect 589398 116651 591448 118972
rect 592028 415428 593928 430800
rect 592028 412948 593928 413528
rect 592028 410578 593928 410898
rect 592028 407872 593928 408528
rect 592028 405502 593928 405822
rect 592028 402872 593928 403452
rect 592028 191683 593928 400972
rect 592028 190294 593928 190983
rect 592028 189082 593928 189804
rect 592028 187870 593928 188592
rect 592028 186658 593928 187380
rect 592028 185446 593928 186168
rect 592028 184234 593928 184956
rect 592028 183022 593928 183744
rect 592028 181810 593928 182532
rect 592028 180598 593928 181320
rect 592028 179386 593928 180108
rect 592028 178174 593928 178896
rect 592028 176962 593928 177684
rect 592028 175750 593928 176472
rect 592028 174538 593928 175260
rect 592028 173326 593928 174048
rect 592028 172114 593928 172836
rect 592028 170902 593928 171624
rect 592028 169239 593928 170412
rect 592028 162928 593928 166291
rect 592028 160807 593928 162227
rect 592028 156721 593928 158898
rect 592028 153517 593928 155259
rect 592028 151127 593928 152562
rect 592028 148819 593928 150098
rect 592028 133428 593928 148119
rect 592028 130948 593928 131528
rect 592028 128578 593928 128898
rect 592028 125872 593928 126528
rect 592028 123502 593928 123822
rect 592028 120872 593928 121452
rect 592028 116651 593928 118972
rect 566228 102748 568128 103328
rect 566228 100378 568128 100698
rect 566228 97672 568128 98328
rect 566228 95302 568128 95622
rect 566228 92672 568128 93252
rect 566228 89056 568128 90772
<< via4 >>
rect 218272 413528 220172 415428
rect 218272 410898 220172 412948
rect 218272 408528 220172 410578
rect 218272 405822 220172 407872
rect 218272 403452 220172 405502
rect 218272 400972 220172 402872
rect 192472 385328 194372 387228
rect 192472 382698 194372 384748
rect 192472 380328 194372 382378
rect 192472 377622 194372 379672
rect 192472 375252 194372 377302
rect 192472 372772 194372 374672
rect 192472 103328 194372 105228
rect 192472 100698 194372 102748
rect 192472 98328 194372 100378
rect 192472 95622 194372 97672
rect 192472 93252 194372 95302
rect 192472 90772 194372 92672
rect 194952 385328 197002 387228
rect 194952 382698 197002 384748
rect 194952 380328 197002 382378
rect 194952 377622 197002 379672
rect 194952 375252 197002 377302
rect 194952 372772 197002 374672
rect 194952 103328 197002 105228
rect 194952 100698 197002 102748
rect 194952 98328 197002 100378
rect 194952 95622 197002 97672
rect 194952 93252 197002 95302
rect 194952 90772 197002 92672
rect 197322 385328 199372 387228
rect 197322 382698 199372 384748
rect 197322 380328 199372 382378
rect 197322 377622 199372 379672
rect 197322 375252 199372 377302
rect 197322 372772 199372 374672
rect 197322 103328 199372 105228
rect 197322 100698 199372 102748
rect 197322 98328 199372 100378
rect 197322 95622 199372 97672
rect 197322 93252 199372 95302
rect 197322 90772 199372 92672
rect 200028 385328 202078 387228
rect 200028 382698 202078 384748
rect 200028 380328 202078 382378
rect 200028 377622 202078 379672
rect 200028 375252 202078 377302
rect 200028 372772 202078 374672
rect 200028 103328 202078 105228
rect 200028 100698 202078 102748
rect 200028 98328 202078 100378
rect 200028 95622 202078 97672
rect 200028 93252 202078 95302
rect 200028 90772 202078 92672
rect 202398 385328 204448 387228
rect 202398 382698 204448 384748
rect 202398 380328 204448 382378
rect 202398 377622 204448 379672
rect 202398 375252 204448 377302
rect 202398 372772 204448 374672
rect 202398 103328 204448 105228
rect 202398 100698 204448 102748
rect 202398 98328 204448 100378
rect 202398 95622 204448 97672
rect 202398 93252 204448 95302
rect 202398 90772 204448 92672
rect 205028 385328 206851 387228
rect 205028 382698 206851 384748
rect 205028 380328 206851 382378
rect 205028 377622 206851 379672
rect 205028 375252 206851 377302
rect 205028 372772 206851 374672
rect 205028 103328 206851 105228
rect 205028 100698 206851 102748
rect 205028 98328 206851 100378
rect 205028 95622 206851 97672
rect 205028 93252 206851 95302
rect 205028 90772 206851 92672
rect 218272 131528 220172 133428
rect 218272 128898 220172 130948
rect 218272 126528 220172 128578
rect 218272 123822 220172 125872
rect 218272 121452 220172 123502
rect 218272 118972 220172 120872
rect 220752 413528 222802 415428
rect 220752 410898 222802 412948
rect 220752 408528 222802 410578
rect 220752 405822 222802 407872
rect 220752 403452 222802 405502
rect 220752 400972 222802 402872
rect 220752 131528 222802 133428
rect 220752 128898 222802 130948
rect 220752 126528 222802 128578
rect 220752 123822 222802 125872
rect 220752 121452 222802 123502
rect 220752 118972 222802 120872
rect 223122 413528 225172 415428
rect 223122 410898 225172 412948
rect 223122 408528 225172 410578
rect 223122 405822 225172 407872
rect 223122 403452 225172 405502
rect 223122 400972 225172 402872
rect 223122 131528 225172 133428
rect 223122 128898 225172 130948
rect 223122 126528 225172 128578
rect 223122 123822 225172 125872
rect 223122 121452 225172 123502
rect 223122 118972 225172 120872
rect 225828 413528 227878 415428
rect 225828 410898 227878 412948
rect 225828 408528 227878 410578
rect 225828 405822 227878 407872
rect 225828 403452 227878 405502
rect 225828 400972 227878 402872
rect 225828 131528 227878 133428
rect 225828 128898 227878 130948
rect 225828 126528 227878 128578
rect 225828 123822 227878 125872
rect 225828 121452 227878 123502
rect 225828 118972 227878 120872
rect 228198 413528 230248 415428
rect 228198 410898 230248 412948
rect 228198 408528 230248 410578
rect 228198 405822 230248 407872
rect 228198 403452 230248 405502
rect 228198 400972 230248 402872
rect 228198 131528 230248 133428
rect 228198 128898 230248 130948
rect 228198 126528 230248 128578
rect 228198 123822 230248 125872
rect 228198 121452 230248 123502
rect 228198 118972 230248 120872
rect 230828 413528 232655 415428
rect 230828 410898 232655 412948
rect 230828 408528 232655 410578
rect 230828 405822 232655 407872
rect 230828 403452 232655 405502
rect 230828 400972 232655 402872
rect 553672 385328 555572 387228
rect 553672 382698 555572 384748
rect 553672 380328 555572 382378
rect 553672 377622 555572 379672
rect 553672 375252 555572 377302
rect 553672 372772 555572 374672
rect 230828 131528 232655 133428
rect 230828 128898 232655 130948
rect 230828 126528 232655 128578
rect 230828 123822 232655 125872
rect 230828 121452 232655 123502
rect 230828 118972 232655 120872
rect 327021 103328 327835 105228
rect 327021 100698 327835 102748
rect 327021 98328 327835 100378
rect 327021 95622 327835 97672
rect 327021 93252 327835 95302
rect 327021 90772 327835 92672
rect 328649 131528 329463 133428
rect 328649 128898 329463 130948
rect 328649 126528 329463 128578
rect 328649 123822 329463 125872
rect 328649 121452 329463 123502
rect 328649 118972 329463 120872
rect 459446 131528 460246 133428
rect 459446 128898 460246 130948
rect 459446 126528 460246 128578
rect 459446 123822 460246 125872
rect 459446 121452 460246 123502
rect 459446 118972 460246 120872
rect 460979 103328 461779 105228
rect 460979 100698 461779 102748
rect 460979 98328 461779 100378
rect 460979 95622 461779 97672
rect 460979 93252 461779 95302
rect 460979 90772 461779 92672
rect 553672 103328 555572 105228
rect 553672 100698 555572 102748
rect 553672 98328 555572 100378
rect 553672 95622 555572 97672
rect 553672 93252 555572 95302
rect 553672 90772 555572 92672
rect 556152 385328 558202 387228
rect 556152 382698 558202 384748
rect 556152 380328 558202 382378
rect 556152 377622 558202 379672
rect 556152 375252 558202 377302
rect 556152 372772 558202 374672
rect 556152 103328 558202 105228
rect 556152 100698 558202 102748
rect 556152 98328 558202 100378
rect 556152 95622 558202 97672
rect 556152 93252 558202 95302
rect 556152 90772 558202 92672
rect 558522 385328 560572 387228
rect 558522 382698 560572 384748
rect 558522 380328 560572 382378
rect 558522 377622 560572 379672
rect 558522 375252 560572 377302
rect 558522 372772 560572 374672
rect 558522 103328 560572 105228
rect 558522 100698 560572 102748
rect 558522 98328 560572 100378
rect 558522 95622 560572 97672
rect 558522 93252 560572 95302
rect 558522 90772 560572 92672
rect 561228 385328 563278 387228
rect 561228 382698 563278 384748
rect 561228 380328 563278 382378
rect 561228 377622 563278 379672
rect 561228 375252 563278 377302
rect 561228 372772 563278 374672
rect 561228 103328 563278 105228
rect 561228 100698 563278 102748
rect 561228 98328 563278 100378
rect 561228 95622 563278 97672
rect 561228 93252 563278 95302
rect 561228 90772 563278 92672
rect 563598 385328 565648 387228
rect 563598 382698 565648 384748
rect 563598 380328 565648 382378
rect 563598 377622 565648 379672
rect 563598 375252 565648 377302
rect 563598 372772 565648 374672
rect 563598 103328 565648 105228
rect 563598 100698 565648 102748
rect 563598 98328 565648 100378
rect 563598 95622 565648 97672
rect 563598 93252 565648 95302
rect 563598 90772 565648 92672
rect 566228 385328 568128 387228
rect 566228 382698 568128 384748
rect 566228 380328 568128 382378
rect 566228 377622 568128 379672
rect 566228 375252 568128 377302
rect 566228 372772 568128 374672
rect 579472 413528 581372 415428
rect 579472 410898 581372 412948
rect 579472 408528 581372 410578
rect 579472 405822 581372 407872
rect 579472 403452 581372 405502
rect 579472 400972 581372 402872
rect 579472 131528 581372 133428
rect 579472 128898 581372 130948
rect 579472 126528 581372 128578
rect 579472 123822 581372 125872
rect 579472 121452 581372 123502
rect 579472 118972 581372 120872
rect 581952 413528 584002 415428
rect 581952 410898 584002 412948
rect 581952 408528 584002 410578
rect 581952 405822 584002 407872
rect 581952 403452 584002 405502
rect 581952 400972 584002 402872
rect 581952 131528 584002 133428
rect 581952 128898 584002 130948
rect 581952 126528 584002 128578
rect 581952 123822 584002 125872
rect 581952 121452 584002 123502
rect 581952 118972 584002 120872
rect 584322 413528 586372 415428
rect 584322 410898 586372 412948
rect 584322 408528 586372 410578
rect 584322 405822 586372 407872
rect 584322 403452 586372 405502
rect 584322 400972 586372 402872
rect 584322 131528 586372 133428
rect 584322 128898 586372 130948
rect 584322 126528 586372 128578
rect 584322 123822 586372 125872
rect 584322 121452 586372 123502
rect 584322 118972 586372 120872
rect 587028 413528 589078 415428
rect 587028 410898 589078 412948
rect 587028 408528 589078 410578
rect 587028 405822 589078 407872
rect 587028 403452 589078 405502
rect 587028 400972 589078 402872
rect 587028 131528 589078 133428
rect 587028 128898 589078 130948
rect 587028 126528 589078 128578
rect 587028 123822 589078 125872
rect 587028 121452 589078 123502
rect 587028 118972 589078 120872
rect 589398 413528 591448 415428
rect 589398 410898 591448 412948
rect 589398 408528 591448 410578
rect 589398 405822 591448 407872
rect 589398 403452 591448 405502
rect 589398 400972 591448 402872
rect 589398 131528 591448 133428
rect 589398 128898 591448 130948
rect 589398 126528 591448 128578
rect 589398 123822 591448 125872
rect 589398 121452 591448 123502
rect 589398 118972 591448 120872
rect 592028 413528 593928 415428
rect 592028 410898 593928 412948
rect 592028 408528 593928 410578
rect 592028 405822 593928 407872
rect 592028 403452 593928 405502
rect 592028 400972 593928 402872
rect 592028 131528 593928 133428
rect 592028 128898 593928 130948
rect 592028 126528 593928 128578
rect 592028 123822 593928 125872
rect 592028 121452 593928 123502
rect 592028 118972 593928 120872
rect 566228 103328 568128 105228
rect 566228 100698 568128 102748
rect 566228 98328 568128 100378
rect 566228 95622 568128 97672
rect 566228 93252 568128 95302
rect 566228 90772 568128 92672
<< metal5 >>
rect 90500 488600 102500 500600
rect 116300 488600 128300 500600
rect 142100 488600 154100 500600
rect 167900 488600 179900 500600
rect 193700 488600 205700 500600
rect 219500 488600 231500 500600
rect 245300 488600 257300 500600
rect 271100 488600 283100 500600
rect 296900 488600 308900 500600
rect 322700 488600 334700 500600
rect 348500 488600 360500 500600
rect 374300 488600 386300 500600
rect 400100 488600 412100 500600
rect 425900 488600 437900 500600
rect 451700 488600 463700 500600
rect 477500 488600 489500 500600
rect 503300 488600 515300 500600
rect 529100 488600 541100 500600
rect 554900 488600 566900 500600
rect 580700 488600 592700 500600
rect 606500 488600 618500 500600
rect 632300 488600 644300 500600
rect 658100 488600 670100 500600
rect 683900 488600 695900 500600
rect 5600 402200 17600 414200
rect 75470 413528 218272 415428
rect 220172 413528 220752 415428
rect 222802 413528 223122 415428
rect 225172 413528 225828 415428
rect 227878 413528 228198 415428
rect 230248 413528 230828 415428
rect 232655 413528 579472 415428
rect 581372 413528 581952 415428
rect 584002 413528 584322 415428
rect 586372 413528 587028 415428
rect 589078 413528 589398 415428
rect 591448 413528 592028 415428
rect 593928 413528 595413 415428
rect 75470 410898 218272 412948
rect 220172 410898 220752 412948
rect 222802 410898 223122 412948
rect 225172 410898 225828 412948
rect 227878 410898 228198 412948
rect 230248 410898 230828 412948
rect 232655 410898 579472 412948
rect 581372 410898 581952 412948
rect 584002 410898 584322 412948
rect 586372 410898 587028 412948
rect 589078 410898 589398 412948
rect 591448 410898 592028 412948
rect 593928 410898 595413 412948
rect 75470 408528 218272 410578
rect 220172 408528 220752 410578
rect 222802 408528 223122 410578
rect 225172 408528 225828 410578
rect 227878 408528 228198 410578
rect 230248 408528 230828 410578
rect 232655 408528 579472 410578
rect 581372 408528 581952 410578
rect 584002 408528 584322 410578
rect 586372 408528 587028 410578
rect 589078 408528 589398 410578
rect 591448 408528 592028 410578
rect 593928 408528 595413 410578
rect 75470 405822 218272 407872
rect 220172 405822 220752 407872
rect 222802 405822 223122 407872
rect 225172 405822 225828 407872
rect 227878 405822 228198 407872
rect 230248 405822 230828 407872
rect 232655 405822 579472 407872
rect 581372 405822 581952 407872
rect 584002 405822 584322 407872
rect 586372 405822 587028 407872
rect 589078 405822 589398 407872
rect 591448 405822 592028 407872
rect 593928 405822 595413 407872
rect 75470 403452 218272 405502
rect 220172 403452 220752 405502
rect 222802 403452 223122 405502
rect 225172 403452 225828 405502
rect 227878 403452 228198 405502
rect 230248 403452 230828 405502
rect 232655 403452 579472 405502
rect 581372 403452 581952 405502
rect 584002 403452 584322 405502
rect 586372 403452 587028 405502
rect 589078 403452 589398 405502
rect 591448 403452 592028 405502
rect 593928 403452 595413 405502
rect 75470 400972 218272 402872
rect 220172 400972 220752 402872
rect 222802 400972 223122 402872
rect 225172 400972 225828 402872
rect 227878 400972 228198 402872
rect 230248 400972 230828 402872
rect 232655 400972 579472 402872
rect 581372 400972 581952 402872
rect 584002 400972 584322 402872
rect 586372 400972 587028 402872
rect 589078 400972 589398 402872
rect 591448 400972 592028 402872
rect 593928 400972 595413 402872
rect 768800 402200 780800 414200
rect 5600 374000 17600 386000
rect 75470 385328 192472 387228
rect 194372 385328 194952 387228
rect 197002 385328 197322 387228
rect 199372 385328 200028 387228
rect 202078 385328 202398 387228
rect 204448 385328 205028 387228
rect 206851 385328 553672 387228
rect 555572 385328 556152 387228
rect 558202 385328 558522 387228
rect 560572 385328 561228 387228
rect 563278 385328 563598 387228
rect 565648 385328 566228 387228
rect 568128 385328 570501 387228
rect 75470 382698 192472 384748
rect 194372 382698 194952 384748
rect 197002 382698 197322 384748
rect 199372 382698 200028 384748
rect 202078 382698 202398 384748
rect 204448 382698 205028 384748
rect 206851 382698 553672 384748
rect 555572 382698 556152 384748
rect 558202 382698 558522 384748
rect 560572 382698 561228 384748
rect 563278 382698 563598 384748
rect 565648 382698 566228 384748
rect 568128 382698 570501 384748
rect 75470 380328 192472 382378
rect 194372 380328 194952 382378
rect 197002 380328 197322 382378
rect 199372 380328 200028 382378
rect 202078 380328 202398 382378
rect 204448 380328 205028 382378
rect 206851 380328 553672 382378
rect 555572 380328 556152 382378
rect 558202 380328 558522 382378
rect 560572 380328 561228 382378
rect 563278 380328 563598 382378
rect 565648 380328 566228 382378
rect 568128 380328 570501 382378
rect 75470 377622 192472 379672
rect 194372 377622 194952 379672
rect 197002 377622 197322 379672
rect 199372 377622 200028 379672
rect 202078 377622 202398 379672
rect 204448 377622 205028 379672
rect 206851 377622 553672 379672
rect 555572 377622 556152 379672
rect 558202 377622 558522 379672
rect 560572 377622 561228 379672
rect 563278 377622 563598 379672
rect 565648 377622 566228 379672
rect 568128 377622 570501 379672
rect 75470 375252 192472 377302
rect 194372 375252 194952 377302
rect 197002 375252 197322 377302
rect 199372 375252 200028 377302
rect 202078 375252 202398 377302
rect 204448 375252 205028 377302
rect 206851 375252 553672 377302
rect 555572 375252 556152 377302
rect 558202 375252 558522 377302
rect 560572 375252 561228 377302
rect 563278 375252 563598 377302
rect 565648 375252 566228 377302
rect 568128 375252 570501 377302
rect 75470 372772 192472 374672
rect 194372 372772 194952 374672
rect 197002 372772 197322 374672
rect 199372 372772 200028 374672
rect 202078 372772 202398 374672
rect 204448 372772 205028 374672
rect 206851 372772 553672 374672
rect 555572 372772 556152 374672
rect 558202 372772 558522 374672
rect 560572 372772 561228 374672
rect 563278 372772 563598 374672
rect 565648 372772 566228 374672
rect 568128 372772 570501 374672
rect 768800 374000 780800 386000
rect 5600 345800 17600 357800
rect 768800 345800 780800 357800
rect 5600 317600 17600 329600
rect 768800 317600 780800 329600
rect 5600 289400 17600 301400
rect 768800 289400 780800 301400
rect 5600 261200 17600 273200
rect 768800 261200 780800 273200
rect 5600 233000 17600 245000
rect 768800 233000 780800 245000
rect 5600 204800 17600 216800
rect 768800 204800 780800 216800
rect 5600 176600 17600 188600
rect 768800 176600 780800 188600
rect 5600 148400 17600 160400
rect 768800 148400 780800 160400
rect 5600 120200 17600 132200
rect 215994 131528 218272 133428
rect 220172 131528 220752 133428
rect 222802 131528 223122 133428
rect 225172 131528 225828 133428
rect 227878 131528 228198 133428
rect 230248 131528 230828 133428
rect 232655 131528 328649 133428
rect 329463 131528 459446 133428
rect 460246 131528 579472 133428
rect 581372 131528 581952 133428
rect 584002 131528 584322 133428
rect 586372 131528 587028 133428
rect 589078 131528 589398 133428
rect 591448 131528 592028 133428
rect 593928 131528 710930 133428
rect 215994 128898 218272 130948
rect 220172 128898 220752 130948
rect 222802 128898 223122 130948
rect 225172 128898 225828 130948
rect 227878 128898 228198 130948
rect 230248 128898 230828 130948
rect 232655 128898 328649 130948
rect 329463 128898 459446 130948
rect 460246 128898 579472 130948
rect 581372 128898 581952 130948
rect 584002 128898 584322 130948
rect 586372 128898 587028 130948
rect 589078 128898 589398 130948
rect 591448 128898 592028 130948
rect 593928 128898 710930 130948
rect 215994 126528 218272 128578
rect 220172 126528 220752 128578
rect 222802 126528 223122 128578
rect 225172 126528 225828 128578
rect 227878 126528 228198 128578
rect 230248 126528 230828 128578
rect 232655 126528 328649 128578
rect 329463 126528 459446 128578
rect 460246 126528 579472 128578
rect 581372 126528 581952 128578
rect 584002 126528 584322 128578
rect 586372 126528 587028 128578
rect 589078 126528 589398 128578
rect 591448 126528 592028 128578
rect 593928 126528 710930 128578
rect 215994 123822 218272 125872
rect 220172 123822 220752 125872
rect 222802 123822 223122 125872
rect 225172 123822 225828 125872
rect 227878 123822 228198 125872
rect 230248 123822 230828 125872
rect 232655 123822 328649 125872
rect 329463 123822 459446 125872
rect 460246 123822 579472 125872
rect 581372 123822 581952 125872
rect 584002 123822 584322 125872
rect 586372 123822 587028 125872
rect 589078 123822 589398 125872
rect 591448 123822 592028 125872
rect 593928 123822 710930 125872
rect 215994 121452 218272 123502
rect 220172 121452 220752 123502
rect 222802 121452 223122 123502
rect 225172 121452 225828 123502
rect 227878 121452 228198 123502
rect 230248 121452 230828 123502
rect 232655 121452 328649 123502
rect 329463 121452 459446 123502
rect 460246 121452 579472 123502
rect 581372 121452 581952 123502
rect 584002 121452 584322 123502
rect 586372 121452 587028 123502
rect 589078 121452 589398 123502
rect 591448 121452 592028 123502
rect 593928 121452 710930 123502
rect 75376 119599 85827 120399
rect 5600 92000 17600 104000
rect 75376 91275 83762 92075
rect 82962 86052 83762 91275
rect 85027 88082 85827 119599
rect 215994 118972 218272 120872
rect 220172 118972 220752 120872
rect 222802 118972 223122 120872
rect 225172 118972 225828 120872
rect 227878 118972 228198 120872
rect 230248 118972 230828 120872
rect 232655 118972 328649 120872
rect 329463 118972 459446 120872
rect 460246 118972 579472 120872
rect 581372 118972 581952 120872
rect 584002 118972 584322 120872
rect 586372 118972 587028 120872
rect 589078 118972 589398 120872
rect 591448 118972 592028 120872
rect 593928 118972 710930 120872
rect 768800 120200 780800 132200
rect 190699 103328 192472 105228
rect 194372 103328 194952 105228
rect 197002 103328 197322 105228
rect 199372 103328 200028 105228
rect 202078 103328 202398 105228
rect 204448 103328 205028 105228
rect 206851 103328 327021 105228
rect 327835 103328 460979 105228
rect 461779 103328 553672 105228
rect 555572 103328 556152 105228
rect 558202 103328 558522 105228
rect 560572 103328 561228 105228
rect 563278 103328 563598 105228
rect 565648 103328 566228 105228
rect 568128 103328 710930 105228
rect 190699 100698 192472 102748
rect 194372 100698 194952 102748
rect 197002 100698 197322 102748
rect 199372 100698 200028 102748
rect 202078 100698 202398 102748
rect 204448 100698 205028 102748
rect 206851 100698 327021 102748
rect 327835 100698 460979 102748
rect 461779 100698 553672 102748
rect 555572 100698 556152 102748
rect 558202 100698 558522 102748
rect 560572 100698 561228 102748
rect 563278 100698 563598 102748
rect 565648 100698 566228 102748
rect 568128 100698 710930 102748
rect 190699 98328 192472 100378
rect 194372 98328 194952 100378
rect 197002 98328 197322 100378
rect 199372 98328 200028 100378
rect 202078 98328 202398 100378
rect 204448 98328 205028 100378
rect 206851 98328 327021 100378
rect 327835 98328 460979 100378
rect 461779 98328 553672 100378
rect 555572 98328 556152 100378
rect 558202 98328 558522 100378
rect 560572 98328 561228 100378
rect 563278 98328 563598 100378
rect 565648 98328 566228 100378
rect 568128 98328 710930 100378
rect 190699 95622 192472 97672
rect 194372 95622 194952 97672
rect 197002 95622 197322 97672
rect 199372 95622 200028 97672
rect 202078 95622 202398 97672
rect 204448 95622 205028 97672
rect 206851 95622 327021 97672
rect 327835 95622 460979 97672
rect 461779 95622 553672 97672
rect 555572 95622 556152 97672
rect 558202 95622 558522 97672
rect 560572 95622 561228 97672
rect 563278 95622 563598 97672
rect 565648 95622 566228 97672
rect 568128 95622 710930 97672
rect 190699 93252 192472 95302
rect 194372 93252 194952 95302
rect 197002 93252 197322 95302
rect 199372 93252 200028 95302
rect 202078 93252 202398 95302
rect 204448 93252 205028 95302
rect 206851 93252 327021 95302
rect 327835 93252 460979 95302
rect 461779 93252 553672 95302
rect 555572 93252 556152 95302
rect 558202 93252 558522 95302
rect 560572 93252 561228 95302
rect 563278 93252 563598 95302
rect 565648 93252 566228 95302
rect 568128 93252 710930 95302
rect 190699 90772 192472 92672
rect 194372 90772 194952 92672
rect 197002 90772 197322 92672
rect 199372 90772 200028 92672
rect 202078 90772 202398 92672
rect 204448 90772 205028 92672
rect 206851 90772 327021 92672
rect 327835 90772 460979 92672
rect 461779 90772 553672 92672
rect 555572 90772 556152 92672
rect 558202 90772 558522 92672
rect 560572 90772 561228 92672
rect 563278 90772 563598 92672
rect 565648 90772 566228 92672
rect 568128 90772 710930 92672
rect 768800 92000 780800 104000
rect 85027 87282 155240 88082
rect 82962 85252 155240 86052
rect 90500 5600 102500 17600
rect 116300 5600 128300 17600
rect 142100 5600 154100 17600
rect 167900 5600 179900 17600
rect 193700 5600 205700 17600
rect 219500 5600 231500 17600
rect 245300 5600 257300 17600
rect 271100 5600 283100 17600
rect 296900 5600 308900 17600
rect 322700 5600 334700 17600
rect 348500 5600 360500 17600
rect 374300 5600 386300 17600
rect 400100 5600 412100 17600
rect 425900 5600 437900 17600
rect 451700 5600 463700 17600
rect 477500 5600 489500 17600
rect 503300 5600 515300 17600
rect 529100 5600 541100 17600
rect 554900 5600 566900 17600
rect 580700 5600 592700 17600
rect 606500 5600 618500 17600
rect 632300 5600 644300 17600
rect 658100 5600 670100 17600
rect 683900 5600 695900 17600
use chip_half_frame  chip_half_frame_0
timestamp 1766089602
transform 1 0 0 0 1 0
box 5200 5200 781200 501000
use copyright_block  copyright_block_0
timestamp 1764012043
transform 1 0 64235 0 1 6580
box 0 570 19550 9198
use gf180mcu_ocd_ip_sram__sram256x8m8wm1  gf180mcu_ocd_ip_sram__sram256x8m8wm1_0 $PDKPATH/libs.ref/gf180mcu_ocd_ip_sram/mag
timestamp 1765987700
transform 1 0 485767 0 1 147257
box 0 0 60260 44986
use gf180mcu_ocd_ip_sram__sram256x8m8wm1  gf180mcu_ocd_ip_sram__sram256x8m8wm1_1
timestamp 1765987700
transform 1 0 601323 0 1 147256
box 0 0 60260 44986
use gf180mcu_ocd_ip_sram__sram512x8m8wm1  gf180mcu_ocd_ip_sram__sram512x8m8wm1_0 $PDKPATH/libs.ref/gf180mcu_ocd_ip_sram/mag
timestamp 1765987700
transform 1 0 245134 0 1 147760
box 0 0 60260 64378
use gf180mcu_ocd_ip_sram__sram1024x8m8wm1  gf180mcu_ocd_ip_sram__sram1024x8m8wm1_0 $PDKPATH/libs.ref/gf180mcu_ocd_ip_sram/mag
timestamp 1765987700
transform 1 0 120566 0 1 147758
box 0 0 60260 103162
use horz_via_program_input  horz_via_program_input_0
timestamp 1765074470
transform 1 0 0 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_2
timestamp 1765074470
transform 1 0 103200 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_3
timestamp 1765074470
transform 1 0 129000 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_4
timestamp 1765074470
transform 1 0 154801 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_5
timestamp 1765074470
transform 1 0 180600 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_6
timestamp 1765074470
transform 1 0 206400 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_7
timestamp 1765074470
transform 1 0 232200 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_8
timestamp 1765074470
transform 1 0 258000 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_9
timestamp 1765074470
transform 1 0 283800 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_10
timestamp 1765074470
transform 1 0 309600 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_11
timestamp 1765074470
transform 1 0 335400 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_12
timestamp 1765074470
transform 1 0 361200 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_13
timestamp 1765074470
transform 1 0 387000 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_14
timestamp 1765074470
transform 1 0 464400 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_15
timestamp 1765074470
transform 1 0 490200 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_16
timestamp 1765074470
transform 1 0 516000 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_17
timestamp 1765074470
transform 1 0 541800 0 1 0
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_18
timestamp 1765074470
transform 1 0 541800 0 -1 506200
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_19
timestamp 1765074470
transform 1 0 516000 0 -1 506200
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_20
timestamp 1765074470
transform 1 0 490200 0 -1 506200
box 141282 75235 154691 75385
use horz_via_program_input  horz_via_program_input_21
timestamp 1765074470
transform 1 0 464400 0 -1 506200
box 141282 75235 154691 75385
use horz_via_program_output  horz_via_program_output_0
timestamp 1765074952
transform 1 0 1 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_1
timestamp 1765074952
transform 1 0 -25799 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_2
timestamp 1765074952
transform 1 0 -51599 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_3
timestamp 1765074952
transform 1 0 -77399 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_4
timestamp 1765074952
transform 1 0 -103199 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_5
timestamp 1765074952
transform 1 0 -128999 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_6
timestamp 1765074952
transform 1 0 -154799 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_7
timestamp 1765074952
transform 1 0 -180599 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_8
timestamp 1765074952
transform 1 0 -206399 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_9
timestamp 1765074952
transform 1 0 -232199 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_10
timestamp 1765074952
transform 1 0 -257999 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_11
timestamp 1765074952
transform 1 0 -283799 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_12
timestamp 1765074952
transform 1 0 -361199 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_13
timestamp 1765074952
transform 1 0 -386999 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_14
timestamp 1765074952
transform 1 0 -412799 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_15
timestamp 1765074952
transform 1 0 -438599 0 1 0
box 528281 430815 541692 430965
use horz_via_program_output  horz_via_program_output_16
timestamp 1765074952
transform 1 0 -361200 0 -1 506200
box 528281 430815 541692 430965
use lvlshift_down  lvlshift_down_0
timestamp 1766090161
transform 0 -1 184611 1 0 81921
box -1221 1570 3231 3370
use ocd_mux_array  ocd_mux_array_0
timestamp 1765233513
transform 1 0 -937 0 1 194
box 467911 148869 484450 151238
use ocd_mux_array  ocd_mux_array_1
timestamp 1765233513
transform 1 0 -158761 0 1 -110
box 467911 148869 484450 151238
use ocd_via2_3x  ocd_via2_3x_0
timestamp 1765059587
transform 1 0 0 0 1 0
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_1
timestamp 1765059587
transform 1 0 64920 0 1 -200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_2
timestamp 1765059587
transform 1 0 -1827 0 1 -9399
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_3
timestamp 1765059587
transform 1 0 168112 0 1 -599
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_4
timestamp 1765059587
transform 1 0 195997 0 1 -800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_5
timestamp 1765059587
transform 1 0 219684 0 1 -1000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_6
timestamp 1765059587
transform 1 0 245513 0 1 -1200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_7
timestamp 1765059587
transform 1 0 271317 0 1 -1400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_8
timestamp 1765059587
transform 1 0 297076 0 1 -1600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_9
timestamp 1765059587
transform 1 0 322886 0 1 -1800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_10
timestamp 1765059587
transform 1 0 348696 0 1 -2000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_11
timestamp 1765059587
transform 1 0 374536 0 1 -2200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_12
timestamp 1765059587
transform 1 0 400315 0 1 -2400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_13
timestamp 1765059587
transform 1 0 426081 0 1 -2600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_14
timestamp 1765059587
transform 1 0 451926 0 1 -2800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_15
timestamp 1765059587
transform 1 0 529324 0 1 -3000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_16
timestamp 1765059587
transform 1 0 556879 0 1 -3200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_17
timestamp 1765059587
transform 1 0 580936 0 1 -3400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_18
timestamp 1765059587
transform 1 0 606743 0 1 -3600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_19
timestamp 1765059587
transform 1 0 607372 0 1 -5400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_20
timestamp 1765059587
transform 1 0 607384 0 1 14644
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_21
timestamp 1765059587
transform 1 0 608075 0 1 -5600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_22
timestamp 1765059587
transform 1 0 608088 0 1 42843
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_23
timestamp 1765059587
transform 1 0 608660 0 1 -5800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_24
timestamp 1765059587
transform 1 0 608684 0 1 71044
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_25
timestamp 1765059587
transform 1 0 609325 0 1 -6000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_26
timestamp 1765059587
transform 1 0 609334 0 1 99244
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_27
timestamp 1765059587
transform 1 0 609745 0 1 -3798
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_28
timestamp 1765059587
transform 1 0 610116 0 1 -4001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_29
timestamp 1765059587
transform 1 0 610446 0 1 -4197
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_30
timestamp 1765059587
transform 1 0 610802 0 1 -4400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_31
timestamp 1765059587
transform 1 0 611162 0 1 -4599
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_32
timestamp 1765059587
transform 1 0 611537 0 1 -4799
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_33
timestamp 1765059587
transform 1 0 611921 0 1 -5000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_34
timestamp 1765059587
transform 1 0 612296 0 1 -5201
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_35
timestamp 1765059587
transform 1 0 612357 0 1 127444
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_36
timestamp 1765059587
transform 1 0 611975 0 1 155644
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_37
timestamp 1765059587
transform 1 0 611589 0 1 183844
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_38
timestamp 1765059587
transform 1 0 611227 0 1 212044
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_39
timestamp 1765059587
transform 1 0 610843 0 1 283649
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_40
timestamp 1765059587
transform 1 0 610465 0 1 283186
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_41
timestamp 1765059587
transform 1 0 610096 0 1 282694
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_42
timestamp 1765059587
transform 1 0 609711 0 1 282282
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_43
timestamp 1765059587
transform 1 0 606770 0 1 283648
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_44
timestamp 1765059587
transform 1 0 580928 0 1 283184
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_45
timestamp 1765059587
transform 1 0 555137 0 1 282695
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_46
timestamp 1765059587
transform 1 0 529375 0 1 282280
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_47
timestamp 1765059587
transform 1 0 393676 0 -1 286763
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_48
timestamp 1765059587
transform 1 0 392599 0 -1 285150
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_49
timestamp 1765059587
transform 1 0 391613 0 -1 286551
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_50
timestamp 1765059587
transform 1 0 389594 0 -1 286353
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_51
timestamp 1765059587
transform 1 0 387582 0 -1 286155
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_52
timestamp 1765059587
transform 1 0 385602 0 -1 285957
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_53
timestamp 1765059587
transform 1 0 383555 0 -1 285755
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_54
timestamp 1765059587
transform 1 0 381485 0 -1 285557
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_55
timestamp 1765059587
transform 1 0 379610 0 -1 285355
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_56
timestamp 1765059587
transform 1 0 390553 0 -1 284944
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_57
timestamp 1765059587
transform 1 0 388568 0 -1 284754
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_58
timestamp 1765059587
transform 1 0 386553 0 -1 284552
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_59
timestamp 1765059587
transform 1 0 384608 0 -1 284354
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_60
timestamp 1765059587
transform 1 0 382581 0 -1 284156
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_61
timestamp 1765059587
transform 1 0 380581 0 -1 283954
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_62
timestamp 1765059587
transform 1 0 378573 0 -1 283756
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_63
timestamp 1765059587
transform 1 0 220762 0 1 -9200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_64
timestamp 1765059587
transform 1 0 222774 0 1 -9001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_65
timestamp 1765059587
transform 1 0 224749 0 1 -8802
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_66
timestamp 1765059587
transform 1 0 226760 0 1 -8601
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_67
timestamp 1765059587
transform 1 0 228765 0 1 -8402
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_68
timestamp 1765059587
transform 1 0 230745 0 1 -8203
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_69
timestamp 1765059587
transform 1 0 232755 0 1 -8005
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_70
timestamp 1765059587
transform 1 0 234725 0 1 -7801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_71
timestamp 1765059587
transform 1 0 223741 0 1 -7400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_72
timestamp 1765059587
transform 1 0 225759 0 1 -7198
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_73
timestamp 1765059587
transform 1 0 227788 0 1 -6999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_74
timestamp 1765059587
transform 1 0 229772 0 1 -6798
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_75
timestamp 1765059587
transform 1 0 231772 0 1 -6600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_76
timestamp 1765059587
transform 1 0 233769 0 1 -6401
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_77
timestamp 1765059587
transform 1 0 235771 0 1 -6199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_78
timestamp 1765059587
transform 1 0 32059 0 1 -3598
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_79
timestamp 1765059587
transform 1 0 32762 0 1 -5196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_80
timestamp 1765059587
transform 1 0 33507 0 1 -7601
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_81
timestamp 1765059587
transform 1 0 38813 0 1 -7400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_82
timestamp 1765059587
transform 1 0 39208 0 1 -3407
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_83
timestamp 1765059587
transform 1 0 39580 0 1 -5000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_84
timestamp 1765059587
transform 1 0 39861 0 1 -4799
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_85
timestamp 1765059587
transform 1 0 40188 0 1 -3198
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_86
timestamp 1765059587
transform 1 0 40618 0 1 -7203
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_87
timestamp 1765059587
transform 1 0 46310 0 1 -6999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_88
timestamp 1765059587
transform 1 0 47086 0 1 -4600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_89
timestamp 1765059587
transform 1 0 47443 0 1 -2999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_90
timestamp 1765059587
transform 1 0 50274 0 1 4
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_91
timestamp 1765059587
transform 1 0 51037 0 1 -401
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_92
timestamp 1765059587
transform 1 0 51482 0 1 -597
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_93
timestamp 1765059587
transform 1 0 52314 0 1 -1600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_94
timestamp 1765059587
transform 1 0 53494 0 1 -1801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_95
timestamp 1765059587
transform 1 0 54706 0 1 -2001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_96
timestamp 1765059587
transform 1 0 59159 0 1 -197
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_97
timestamp 1765059587
transform 1 0 65991 0 1 -5401
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_98
timestamp 1765059587
transform 1 0 68366 0 1 -800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_99
timestamp 1765059587
transform 1 0 68843 0 1 -1003
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_100
timestamp 1765059587
transform 1 0 69345 0 1 -1199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_101
timestamp 1765059587
transform 1 0 70114 0 1 -1397
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_102
timestamp 1765059587
transform 1 0 73555 0 1 -2802
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_103
timestamp 1765059587
transform 1 0 74032 0 1 -4398
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_104
timestamp 1765059587
transform 1 0 74593 0 1 -6805
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_105
timestamp 1765059587
transform 1 0 80105 0 1 -6603
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_106
timestamp 1765059587
transform 1 0 80551 0 1 -2600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_107
timestamp 1765059587
transform 1 0 80912 0 1 -4199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_108
timestamp 1765059587
transform 1 0 81343 0 1 -4001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_109
timestamp 1765059587
transform 1 0 81712 0 1 -2400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_110
timestamp 1765059587
transform 1 0 82126 0 1 -6400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_111
timestamp 1765059587
transform 1 0 87850 0 1 -6201
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_112
timestamp 1765059587
transform 1 0 88421 0 1 -3800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_113
timestamp 1765059587
transform 1 0 88912 0 1 -2196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_114
timestamp 1765059587
transform 1 0 212986 0 1 -3800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_115
timestamp 1765059587
transform 1 0 213477 0 1 -2196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_116
timestamp 1765059587
transform 1 0 206277 0 1 -2400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_117
timestamp 1765059587
transform 1 0 205908 0 1 -4001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_118
timestamp 1765059587
transform 1 0 205477 0 1 -4199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_119
timestamp 1765059587
transform 1 0 205116 0 1 -2600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_120
timestamp 1765059587
transform 1 0 198597 0 1 -4398
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_121
timestamp 1765059587
transform 1 0 198120 0 1 -2802
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_122
timestamp 1765059587
transform 1 0 194679 0 1 -1397
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_123
timestamp 1765059587
transform 1 0 193910 0 1 -1199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_124
timestamp 1765059587
transform 1 0 193408 0 1 -1003
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_125
timestamp 1765059587
transform 1 0 192931 0 1 -800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_126
timestamp 1765059587
transform 1 0 178059 0 1 -1801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_127
timestamp 1765059587
transform 1 0 179271 0 1 -2001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_128
timestamp 1765059587
transform 1 0 183724 0 1 -197
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_129
timestamp 1765059587
transform 1 0 172008 0 1 -2999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_130
timestamp 1765059587
transform 1 0 174839 0 1 4
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_131
timestamp 1765059587
transform 1 0 175602 0 1 -401
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_132
timestamp 1765059587
transform 1 0 176047 0 1 -597
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_133
timestamp 1765059587
transform 1 0 176879 0 1 -1600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_134
timestamp 1765059587
transform 1 0 163773 0 1 -3407
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_135
timestamp 1765059587
transform 1 0 164753 0 1 -3198
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_136
timestamp 1765059587
transform 1 0 156624 0 1 -3598
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_137
timestamp 1765059587
transform 1 0 212415 0 1 -7801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_138
timestamp 1765059587
transform 1 0 206691 0 1 -8000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_139
timestamp 1765059587
transform 1 0 199158 0 1 -8405
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_140
timestamp 1765059587
transform 1 0 204670 0 1 -8203
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_141
timestamp 1765059587
transform 1 0 190556 0 1 -5601
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_142
timestamp 1765059587
transform 1 0 170875 0 1 -8599
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_143
timestamp 1765059587
transform 1 0 171651 0 1 -4600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_144
timestamp 1765059587
transform 1 0 163378 0 1 -9000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_145
timestamp 1765059587
transform 1 0 164145 0 1 -5000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_146
timestamp 1765059587
transform 1 0 164426 0 1 -4799
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_147
timestamp 1765059587
transform 1 0 165183 0 1 -8803
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_148
timestamp 1765059587
transform 1 0 157327 0 1 -5196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_149
timestamp 1765059587
transform 1 0 158072 0 1 -9201
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_150
timestamp 1765059587
transform 1 0 397259 0 1 -3598
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_151
timestamp 1765059587
transform 1 0 397962 0 1 -5196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_152
timestamp 1765059587
transform 1 0 398707 0 1 -7601
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_153
timestamp 1765059587
transform 1 0 404408 0 1 -3407
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_154
timestamp 1765059587
transform 1 0 405388 0 1 -3198
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_155
timestamp 1765059587
transform 1 0 404013 0 1 -7400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_156
timestamp 1765059587
transform 1 0 404780 0 1 -5000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_157
timestamp 1765059587
transform 1 0 405061 0 1 -4799
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_158
timestamp 1765059587
transform 1 0 405818 0 1 -7203
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_159
timestamp 1765059587
transform 1 0 412643 0 1 -2999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_160
timestamp 1765059587
transform 1 0 411510 0 1 -6999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_161
timestamp 1765059587
transform 1 0 412286 0 1 -4600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_162
timestamp 1765059587
transform 1 0 431191 0 1 -5801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_163
timestamp 1765059587
transform 1 0 439232 0 1 -4398
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_164
timestamp 1765059587
transform 1 0 438755 0 1 -2802
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_165
timestamp 1765059587
transform 1 0 439793 0 1 -6805
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_166
timestamp 1765059587
transform 1 0 445305 0 1 -6603
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_167
timestamp 1765059587
transform 1 0 446543 0 1 -4001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_168
timestamp 1765059587
transform 1 0 446112 0 1 -4199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_169
timestamp 1765059587
transform 1 0 447326 0 1 -6400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_170
timestamp 1765059587
transform 1 0 453621 0 1 -3800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_171
timestamp 1765059587
transform 1 0 453050 0 1 -6201
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_172
timestamp 1765059587
transform 1 0 415474 0 1 4
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_173
timestamp 1765059587
transform 1 0 569668 0 1 -2196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_174
timestamp 1765059587
transform 1 0 416682 0 1 -597
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_175
timestamp 1765059587
transform 1 0 417514 0 1 -1600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_176
timestamp 1765059587
transform 1 0 418694 0 1 -1801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_177
timestamp 1765059587
transform 1 0 419906 0 1 -2001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_178
timestamp 1765059587
transform 1 0 424359 0 1 -197
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_179
timestamp 1765059587
transform 1 0 435314 0 1 -1397
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_180
timestamp 1765059587
transform 1 0 434545 0 1 -1199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_181
timestamp 1765059587
transform 1 0 434043 0 1 -1003
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_182
timestamp 1765059587
transform 1 0 433566 0 1 -800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_183
timestamp 1765059587
transform 1 0 446912 0 1 -2400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_184
timestamp 1765059587
transform 1 0 445751 0 1 -2600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_185
timestamp 1765059587
transform 1 0 454112 0 1 -2196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_186
timestamp 1765059587
transform 1 0 569177 0 1 -3800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_187
timestamp 1765059587
transform 1 0 561307 0 1 -2600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_188
timestamp 1765059587
transform 1 0 561668 0 1 -4199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_189
timestamp 1765059587
transform 1 0 562099 0 1 -4001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_190
timestamp 1765059587
transform 1 0 562468 0 1 -2400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_191
timestamp 1765059587
transform 1 0 554311 0 1 -2802
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_192
timestamp 1765059587
transform 1 0 554788 0 1 -4398
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_193
timestamp 1765059587
transform 1 0 546747 0 1 -6001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_194
timestamp 1765059587
transform 1 0 549122 0 1 -800
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_195
timestamp 1765059587
transform 1 0 549599 0 1 -1003
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_196
timestamp 1765059587
transform 1 0 550101 0 1 -1199
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_197
timestamp 1765059587
transform 1 0 550870 0 1 -1397
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_198
timestamp 1765059587
transform 1 0 539915 0 1 -197
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_199
timestamp 1765059587
transform 1 0 534250 0 1 -1801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_200
timestamp 1765059587
transform 1 0 533070 0 1 -1600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_201
timestamp 1765059587
transform 1 0 532238 0 1 -597
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_202
timestamp 1765059587
transform 1 0 221762 0 1 -7600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_203
timestamp 1765059587
transform 1 0 531030 0 1 4
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_204
timestamp 1765059587
transform 1 0 535462 0 1 -2001
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_205
timestamp 1765059587
transform 1 0 528199 0 1 -2999
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_206
timestamp 1765059587
transform 1 0 527842 0 1 -4600
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_207
timestamp 1765059587
transform 1 0 520336 0 1 -5000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_208
timestamp 1765059587
transform 1 0 520944 0 1 -3198
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_209
timestamp 1765059587
transform 1 0 519964 0 1 -3407
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_210
timestamp 1765059587
transform 1 0 520617 0 1 -4799
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_211
timestamp 1765059587
transform 1 0 513518 0 1 -5196
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_212
timestamp 1765059587
transform 1 0 512815 0 1 -3598
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_213
timestamp 1765059587
transform 1 0 562882 0 1 -8000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_214
timestamp 1765059587
transform 1 0 568606 0 1 -7801
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_215
timestamp 1765059587
transform 1 0 555349 0 1 -8405
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_216
timestamp 1765059587
transform 1 0 560861 0 1 -8203
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_217
timestamp 1765059587
transform 1 0 527066 0 1 -8599
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_218
timestamp 1765059587
transform 1 0 519569 0 1 -9000
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_219
timestamp 1765059587
transform 1 0 521374 0 1 -8803
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_220
timestamp 1765059587
transform 1 0 514263 0 1 -9201
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_221
timestamp 1765059587
transform 1 0 218412 0 1 -9400
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_222
timestamp 1765059587
transform 1 0 376008 0 -1 283355
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_223
timestamp 1765059587
transform 1 0 376057 0 1 4033
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_224
timestamp 1765059587
transform 1 0 -2207 0 1 -9599
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_225
timestamp 1765059587
transform 1 0 -2391 0 1 29412
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_226
timestamp 1765059587
transform 1 0 -1996 0 1 85814
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_227
timestamp 1765059587
transform 1 0 50669 0 1 200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_228
timestamp 1765059587
transform 1 0 -732 0 1 200
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_229
timestamp 1765059587
transform 1 0 -922 0 1 57612
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_230
timestamp 1765059587
transform 1 0 218399 0 1 3716
box 89752 146428 90065 146528
use simple_por  simple_por_0 ../ip/simple_por/mag
timestamp 1766089602
transform 1 0 155176 0 1 79368
box 0 0 25156 8716
use vert_via_program_input  vert_via_program_input_0
timestamp 1765074735
transform 1 0 0 0 1 0
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_1
timestamp 1765074735
transform 1 0 0 0 1 28200
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_2
timestamp 1765074735
transform 1 0 0 0 1 56400
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_3
timestamp 1765074735
transform 1 0 0 0 1 84600
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_4
timestamp 1765074735
transform 1 0 0 0 1 112800
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_5
timestamp 1765074735
transform 1 0 0 0 1 141000
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_6
timestamp 1765074735
transform 1 0 0 0 1 169200
box 710929 147580 711109 160994
use vert_via_program_input  vert_via_program_input_7
timestamp 1765074735
transform 1 0 0 0 1 197400
box 710929 147580 711109 160994
<< labels >>
flabel metal4 218408 137047 220108 141487 0 FreeSans 16000 90 0 0 VDD
flabel metal4 192533 137156 194168 141852 0 FreeSans 16000 90 0 0 VSS
flabel metal4 553940 136097 555264 140400 0 FreeSans 16000 90 0 0 VSS
flabel metal4 579591 136097 580915 140400 0 FreeSans 16000 90 0 0 VDD
flabel metal3 120657 141282 120657 141282 0 FreeSans 480 0 0 0 WEN0
flabel metal3 120667 141478 120667 141478 0 FreeSans 480 0 0 0 WEN1
flabel metal3 120677 141676 120677 141676 0 FreeSans 480 0 0 0 WEN2
flabel metal3 120685 141876 120685 141876 0 FreeSans 480 0 0 0 WEN3
flabel metal3 120697 142075 120697 142075 0 FreeSans 480 0 0 0 WEN4
flabel metal3 120694 142278 120694 142278 0 FreeSans 480 0 0 0 WEN5
flabel metal3 120680 142478 120680 142478 0 FreeSans 480 0 0 0 WEN6
flabel metal3 120694 142684 120694 142684 0 FreeSans 480 0 0 0 WEN7
flabel metal3 120670 142874 120670 142874 0 FreeSans 480 0 0 0 D0
flabel metal3 120670 143077 120670 143077 0 FreeSans 480 0 0 0 D1
flabel metal3 120667 143268 120667 143268 0 FreeSans 480 0 0 0 D2
flabel metal3 120665 143471 120665 143471 0 FreeSans 480 0 0 0 D3
flabel metal3 120667 143666 120667 143666 0 FreeSans 480 0 0 0 D4
flabel metal3 120667 143872 120667 143872 0 FreeSans 480 0 0 0 D5
flabel metal3 120655 144072 120655 144072 0 FreeSans 480 0 0 0 D6
flabel metal3 120652 144278 120652 144278 0 FreeSans 480 0 0 0 D7
flabel metal3 120667 144476 120667 144476 0 FreeSans 480 0 0 0 A0
flabel metal3 120665 144674 120665 144674 0 FreeSans 480 0 0 0 A1
flabel metal3 120662 144872 120662 144872 0 FreeSans 480 0 0 0 A2
flabel metal3 120652 145078 120652 145078 0 FreeSans 480 0 0 0 A3
flabel metal3 120652 145276 120652 145276 0 FreeSans 480 0 0 0 A4
flabel metal3 120652 145479 120652 145479 0 FreeSans 480 0 0 0 A5
flabel metal3 120667 145674 120667 145674 0 FreeSans 480 0 0 0 A6
flabel metal3 120655 145877 120655 145877 0 FreeSans 480 0 0 0 A7
flabel metal3 120652 146073 120652 146073 0 FreeSans 480 0 0 0 A8
flabel metal3 120640 146278 120640 146278 0 FreeSans 480 0 0 0 GWEN
flabel metal3 120625 146485 120625 146485 0 FreeSans 480 0 0 0 CLK
flabel metal3 120655 140282 120655 140282 0 FreeSans 480 0 0 0 Q7_512_1
flabel metal3 120669 140076 120669 140076 0 FreeSans 480 0 0 0 Q6_512_1
flabel metal3 120671 139874 120671 139874 0 FreeSans 480 0 0 0 Q5_512_1
flabel metal3 120671 139668 120671 139668 0 FreeSans 480 0 0 0 Q4_512_1
flabel metal3 120644 139472 120644 139472 0 FreeSans 480 0 0 0 Q3_512_1
flabel metal3 120638 139274 120638 139274 0 FreeSans 480 0 0 0 Q2_512_1
flabel metal3 120629 139080 120629 139080 0 FreeSans 480 0 0 0 Q1_512_1
flabel metal3 120653 138878 120653 138878 0 FreeSans 480 0 0 0 Q0_512_1
flabel metal3 467224 137481 467224 137481 0 FreeSans 480 0 0 0 Q1_256_2
flabel metal3 467228 137681 467228 137681 0 FreeSans 480 0 0 0 Q2_256_2
flabel metal3 467245 137875 467245 137875 0 FreeSans 480 0 0 0 Q3_256_2
flabel metal3 467235 138676 467235 138676 0 FreeSans 480 0 0 0 Q7_256_2
flabel metal3 467241 138879 467241 138879 0 FreeSans 480 0 0 0 Q0_256_1
flabel metal3 467235 139074 467235 139074 0 FreeSans 480 0 0 0 Q1_256_1
flabel metal3 467228 139276 467228 139276 0 FreeSans 480 0 0 0 Q2_256_1
flabel metal3 467235 139477 467235 139477 0 FreeSans 480 0 0 0 Q3_256_1
flabel metal3 467216 139879 467216 139879 0 FreeSans 480 0 0 0 Q5_256_1
flabel metal3 467239 140078 467239 140078 0 FreeSans 480 0 0 0 Q6_256_1
flabel metal3 467211 140281 467211 140281 0 FreeSans 480 0 0 0 Q7_256_1
flabel metal3 120684 137078 120684 137078 0 FreeSans 480 0 0 0 select_512
flabel metal3 120707 136873 120707 136873 0 FreeSans 480 0 0 0 select_256
flabel metal3 467223 139683 467223 139683 0 FreeSans 480 0 0 0 Q4_256_1
flabel metal3 467230 138477 467230 138477 0 FreeSans 480 0 0 0 Q6_256_2
flabel metal3 467236 138269 467236 138269 0 FreeSans 480 0 0 0 Q5_256_2
flabel metal3 467251 138074 467251 138074 0 FreeSans 480 0 0 0 Q4_256_2
flabel metal3 467227 137278 467227 137278 0 FreeSans 480 0 0 0 Q0_256_2
flabel metal3 245905 138681 245905 138681 0 FreeSans 480 0 0 0 Q7_512_2
flabel metal3 245907 138478 245907 138478 0 FreeSans 480 0 0 0 Q6_512_2
flabel metal3 245909 138278 245909 138278 0 FreeSans 480 0 0 0 Q5_512_2
flabel metal3 245890 138074 245890 138074 0 FreeSans 480 0 0 0 Q4_512_2
flabel metal3 245899 137879 245899 137879 0 FreeSans 480 0 0 0 Q3_512_2
flabel metal3 245897 137674 245897 137674 0 FreeSans 480 0 0 0 Q2_512_2
flabel metal3 245871 137476 245871 137476 0 FreeSans 480 0 0 0 Q1_512_2
flabel metal3 245857 137283 245857 137283 0 FreeSans 480 0 0 0 Q0_512_2
flabel metal3 155240 141077 155240 141077 0 FreeSans 480 0 0 0 ENA_512_1
flabel metal3 279872 140879 279872 140879 0 FreeSans 480 0 0 0 ENA_512_2
flabel metal3 520480 140671 520480 140671 0 FreeSans 480 0 0 0 ENA_256_1
flabel metal3 636077 140468 636077 140468 0 FreeSans 480 0 0 0 ENA_256_2
flabel metal5 90500 5600 102500 17600 0 FreeSans 24000 0 0 0 clk_PAD
port 1 nsew
flabel metal5 116300 5600 128300 17600 0 FreeSans 24000 0 0 0 rst_n_PAD
port 2 nsew
flabel metal5 142100 5600 154100 17600 0 FreeSans 24000 0 0 0 bidir_PAD[0]
port 3 nsew
flabel metal5 167900 5600 179900 17600 0 FreeSans 24000 0 0 0 bidir_PAD[1]
port 4 ne
flabel metal5 193700 5600 205700 17600 0 FreeSans 24000 0 0 0 VSS
port 5 nsew
flabel metal5 219500 5600 231500 17600 0 FreeSans 24000 0 0 0 VDD
port 6 nsew
flabel metal5 245300 5600 257300 17600 0 FreeSans 24000 0 0 0 bidir_PAD[2]
port 7 nsew
flabel metal5 271100 5600 283100 17600 0 FreeSans 24000 0 0 0 bidir_PAD[3]
port 8 nsew
flabel metal5 296900 5600 308900 17600 0 FreeSans 24000 0 0 0 bidir_PAD[4]
port 9 nsew
flabel metal5 322700 5600 334700 17600 0 FreeSans 24000 0 0 0 bidir_PAD[5]
port 10 nsew
flabel metal5 348500 5600 360500 17600 0 FreeSans 24000 0 0 0 bidir_PAD[6]
port 11 nsew
flabel metal5 374300 5600 386300 17600 0 FreeSans 24000 0 0 0 bidir_PAD[7]
port 12 nsew
flabel metal5 400100 5600 412100 17600 0 FreeSans 24000 0 0 0 bidir_PAD[8]
port 13 nsew
flabel metal5 425900 5600 437900 17600 0 FreeSans 24000 0 0 0 bidir_PAD[9]
port 14 nsew
flabel metal5 451700 5600 463700 17600 0 FreeSans 24000 0 0 0 bidir_PAD[10]
port 15 nsew
flabel metal5 477500 5600 489500 17600 0 FreeSans 24000 0 0 0 bidir_PAD[11]
port 16 nsew
flabel metal5 503300 5600 515300 17600 0 FreeSans 24000 0 0 0 bidir_PAD[12]
port 17 nsew
flabel metal5 529100 5600 541100 17600 0 FreeSans 24000 0 0 0 bidir_PAD[13]
port 18 nsew
flabel metal5 554900 5600 566900 17600 0 FreeSans 24000 0 0 0 DVSS
port 23 nsew
flabel metal5 580700 5600 592700 17600 0 FreeSans 24000 0 0 0 DVDD
port 24 nsew
flabel metal5 606500 5600 618500 17600 0 FreeSans 24000 0 0 0 bidir_PAD[14]
port 25 nsew
flabel metal5 632300 5600 644300 17600 0 FreeSans 24000 0 0 0 bidir_PAD[15]
port 26 nsew
flabel metal5 658100 5600 670100 17600 0 FreeSans 24000 0 0 0 bidir_PAD[16]
port 27 nsew
flabel metal5 683900 5600 695900 17600 0 FreeSans 24000 0 0 0 bidir_PAD[17]
port 28 nsew
flabel metal5 768800 148400 780800 160400 0 FreeSans 24000 0 0 0 bidir_PAD[18]
port 29 nsew
flabel metal5 768800 176600 780800 188600 0 FreeSans 24000 0 0 0 bidir_PAD[19]
port 30 nsew
flabel metal5 768800 204800 780800 216800 0 FreeSans 24000 0 0 0 bidir_PAD[20]
port 31 nsew
flabel metal5 768800 233000 780800 245000 0 FreeSans 24000 0 0 0 bidir_PAD[21]
port 32 nsew
flabel metal5 768800 261200 780800 273200 0 FreeSans 24000 0 0 0 bidir_PAD[22]
port 33 nsew
flabel metal5 768800 289400 780800 301400 0 FreeSans 24000 0 0 0 bidir_PAD[23]
port 34 nsew
flabel metal5 768800 317600 780800 329600 0 FreeSans 24000 0 0 0 bidir_PAD[24]
port 35 nsew
flabel metal5 768800 345800 780800 357800 0 FreeSans 24000 0 0 0 bidir_PAD[25]
port 36 nsew
flabel metal5 683900 488600 695900 500600 0 FreeSans 24000 0 0 0 bidir_PAD[26]
port 37 nsew
flabel metal5 658100 488600 670100 500600 0 FreeSans 24000 0 0 0 bidir_PAD[27]
port 38 nsew
flabel metal5 632300 488600 644300 500600 0 FreeSans 24000 0 0 0 bidir_PAD[28]
port 39 nsew
flabel metal5 606500 488600 618500 500600 0 FreeSans 24000 0 0 0 bidir_PAD[29]
port 40 nsew
flabel metal5 529100 488600 541100 500600 0 FreeSans 24000 0 0 0 bidir_PAD[30]
port 41 nsew
flabel metal5 503300 488600 515300 500600 0 FreeSans 24000 0 0 0 bidir_PAD[31]
port 42 nsew
flabel metal5 477500 488600 489500 500600 0 FreeSans 24000 0 0 0 bidir_PAD[32]
port 43 nsew
flabel metal5 451700 488600 463700 500600 0 FreeSans 24000 0 0 0 bidir_PAD[33]
port 44 nsew
flabel metal5 425900 488600 437900 500600 0 FreeSans 24000 0 0 0 bidir_PAD[34]
port 45 nsew
flabel metal5 400100 488600 412100 500600 0 FreeSans 24000 0 0 0 bidir_PAD[35]
port 46 nsew
flabel metal5 374300 488600 386300 500600 0 FreeSans 24000 0 0 0 bidir_PAD[36]
port 47 nsew
flabel metal5 348500 488600 360500 500600 0 FreeSans 24000 0 0 0 bidir_PAD[37]
port 48 nsew
flabel metal5 322700 488600 334700 500600 0 FreeSans 24000 0 0 0 bidir_PAD[38]
port 49 nsew
flabel metal5 296900 488600 308900 500600 0 FreeSans 24000 0 0 0 bidir_PAD[39]
port 50 nsew
flabel metal5 271100 488600 283100 500600 0 FreeSans 24000 0 0 0 bidir_PAD[40]
port 51 nsew
flabel metal5 245300 488600 257300 500600 0 FreeSans 24000 0 0 0 bidir_PAD[41]
port 52 nsew
flabel metal5 167900 488600 179900 500600 0 FreeSans 24000 0 0 0 bidir_PAD[42]
port 53 nsew
flabel metal5 142100 488600 154100 500600 0 FreeSans 24000 0 0 0 bidir_PAD[43]
port 54 nsew
flabel metal5 116300 488600 128300 500600 0 FreeSans 24000 0 0 0 bidir_PAD[44]
port 55 nsew
flabel metal5 90500 488600 102500 500600 0 FreeSans 24000 0 0 0 bidir_PAD[45]
port 56 nsew
flabel metal5 5600 345800 17600 357800 0 FreeSans 24000 0 0 0 analog_PAD[0]
port 57 nsew
flabel metal5 5600 317600 17600 329600 0 FreeSans 24000 0 0 0 analog_PAD[1]
port 58 nsew
flabel metal5 5600 289400 17600 301400 0 FreeSans 24000 0 0 0 analog_PAD[2]
port 59 nsew
flabel metal5 5600 261200 17600 273200 0 FreeSans 24000 0 0 0 analog_PAD[3]
port 60 nsew
flabel metal5 5600 233000 17600 245000 0 FreeSans 24000 0 0 0 input_PAD[0]
port 61 nsew
flabel metal5 5600 204800 17600 216800 0 FreeSans 24000 0 0 0 input_PAD[1]
port 62 nsew
flabel metal5 5600 176600 17600 188600 0 FreeSans 24000 0 0 0 input_PAD[2]
port 63 nsew
flabel metal5 5600 148400 17600 160400 0 FreeSans 24000 0 0 0 input_PAD[3]
port 64 nsew
flabel metal5 5600 120200 17600 132200 0 FreeSans 24000 0 0 0 DVDD
port 24 nsew
flabel metal5 5600 92000 17600 104000 0 FreeSans 24000 0 0 0 DVSS
port 23 nsew
flabel metal5 5600 402200 17600 414200 0 FreeSans 24000 0 0 0 VDD
port 6 nsew
flabel metal5 5600 374000 17600 386000 0 FreeSans 24000 0 0 0 VSS
port 5 nsew
flabel metal5 219500 488600 231500 500600 0 FreeSans 24000 0 0 0 DVDD
port 24 nsew
flabel metal5 193700 488600 205700 500600 0 FreeSans 24000 0 0 0 DVSS
port 23 nsew
flabel metal5 580700 488600 592700 500600 0 FreeSans 24000 0 0 0 VDD
port 6 nsew
flabel metal5 554900 488600 566900 500600 0 FreeSans 24000 0 0 0 VSS
port 5 nsew
flabel metal5 768800 92000 780800 104000 0 FreeSans 24000 0 0 0 VSS
port 5 nsew
flabel metal5 768800 120200 780800 132200 0 FreeSans 24000 0 0 0 VDD
port 6 nsew
flabel metal5 768800 374000 780800 386000 0 FreeSans 24000 0 0 0 DVSS
port 23 nsew
flabel metal5 768800 402200 780800 414200 0 FreeSans 24000 0 0 0 DVDD
port 24 nsew
<< end >>
