magic
tech gf180mcuD
magscale 1 10
timestamp 1764982451
<< metal2 >>
rect 0 14444 270 14456
rect 0 12568 2 14444
rect 269 12568 270 14444
rect 0 12556 270 12568
rect 0 11964 270 11976
rect 0 9938 2 11964
rect 269 9938 270 11964
rect 0 9926 270 9938
rect 0 9594 270 9606
rect 0 7568 2 9594
rect 269 7568 270 9594
rect 0 7556 270 7568
rect 0 6888 270 6900
rect 0 4862 2 6888
rect 269 4862 270 6888
rect 0 4850 270 4862
rect 0 4518 270 4530
rect 0 2492 2 4518
rect 269 2492 270 4518
rect 0 2480 270 2492
rect 0 1888 270 1900
rect 0 12 2 1888
rect 269 12 270 1888
rect 0 0 270 12
<< via2 >>
rect 2 12568 269 14444
rect 2 9938 269 11964
rect 2 7568 269 9594
rect 2 4862 269 6888
rect 2 2492 269 4518
rect 2 12 269 1888
<< metal3 >>
rect 0 14444 270 14456
rect 0 12568 2 14444
rect 269 12568 270 14444
rect 0 11964 270 12568
rect 0 9938 2 11964
rect 269 9938 270 11964
rect 0 9594 270 9938
rect 0 7568 2 9594
rect 269 7568 270 9594
rect 0 6888 270 7568
rect 0 4862 2 6888
rect 269 4862 270 6888
rect 0 4518 270 4862
rect 0 2492 2 4518
rect 269 2492 270 4518
rect 0 1888 270 2492
rect 0 12 2 1888
rect 269 12 270 1888
rect 0 0 270 12
<< via3 >>
rect 2 12568 269 14444
rect 2 9938 269 11964
rect 2 7568 269 9594
rect 2 4862 269 6888
rect 2 2492 269 4518
rect 2 12 269 1888
<< metal4 >>
rect 0 14444 270 14456
rect 0 12568 2 14444
rect 269 12568 270 14444
rect 0 12556 270 12568
rect 0 11964 270 11976
rect 0 9938 2 11964
rect 269 9938 270 11964
rect 0 9926 270 9938
rect 0 9594 270 9606
rect 0 7568 2 9594
rect 269 7568 270 9594
rect 0 7556 270 7568
rect 0 6888 270 6900
rect 0 4862 2 6888
rect 269 4862 270 6888
rect 0 4850 270 4862
rect 0 4518 270 4530
rect 0 2492 2 4518
rect 269 2492 270 4518
rect 0 2480 270 2492
rect 0 1888 270 1900
rect 0 12 2 1888
rect 269 12 270 1888
rect 0 0 270 12
<< via4 >>
rect 2 12568 268 14444
rect 2 9938 268 11964
rect 2 7568 268 9594
rect 2 4862 268 6888
rect 2 2492 268 4518
rect 2 12 268 1888
<< metal5 >>
rect 0 14444 270 14456
rect 0 12568 2 14444
rect 268 12568 270 14444
rect 0 12556 270 12568
rect 0 11964 270 11976
rect 0 9938 2 11964
rect 268 9938 270 11964
rect 0 9926 270 9938
rect 0 9594 270 9606
rect 0 7568 2 9594
rect 268 7568 270 9594
rect 0 7556 270 7568
rect 0 6888 270 6900
rect 0 4862 2 6888
rect 268 4862 270 6888
rect 0 4850 270 4862
rect 0 4518 270 4530
rect 0 2492 2 4518
rect 268 2492 270 4518
rect 0 2480 270 2492
rect 0 1888 270 1900
rect 0 12 2 1888
rect 268 12 270 1888
rect 0 0 270 12
<< properties >>
string flatten true
<< end >>
