magic
tech gf180mcuD
magscale 1 10
timestamp 1765317384
<< checkpaint >>
rect -2000 -2000 788400 508200
<< psubdiff >>
tri 0 504400 1800 506200 se
rect 1800 504400 784600 506200
tri 784600 504400 786400 506200 sw
rect 0 503000 786400 504400
rect 0 3200 3200 503000
rect 783200 3200 786400 503000
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal1 >>
tri 939 505339 1800 506200 se
rect 1800 505339 784600 506200
tri 665 505065 939 505339 se
rect 939 505065 784600 505339
tri 619 505019 665 505065 se
rect 665 505019 784600 505065
tri 299 504699 619 505019 se
rect 619 504699 784600 505019
tri 0 504400 299 504699 se
rect 299 504400 784600 504699
tri 784600 504400 786400 506200 sw
rect 0 503200 786400 504400
rect 0 3000 3000 503200
tri 3000 503000 3200 503200 nw
tri 783200 503000 783400 503200 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 503200
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal2 >>
tri 1288 505688 1800 506200 se
rect 1800 505688 784600 506200
tri 928 505328 1288 505688 se
rect 1288 505328 784600 505688
tri 568 504968 928 505328 se
rect 928 504968 784600 505328
tri 0 504400 568 504968 se
rect 568 504400 784600 504968
tri 784600 504400 786400 506200 sw
rect 0 503000 786400 504400
rect 0 3200 3200 503000
rect 783200 3200 786400 503000
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal3 >>
tri 0 504400 1800 506200 se
rect 1800 504400 784600 506200
tri 784600 504400 786400 506200 sw
rect 0 503200 786400 504400
rect 0 3000 3000 503200
tri 3000 503000 3200 503200 nw
tri 783200 503000 783400 503200 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 503200
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal4 >>
tri 0 504400 1800 506200 se
rect 1800 504400 784600 506200
tri 784600 504400 786400 506200 sw
rect 0 503000 786400 504400
rect 0 3200 3200 503000
rect 783200 3200 786400 503000
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal5 >>
tri 0 504400 1800 506200 se
rect 1800 504400 784600 506200
tri 784600 504400 786400 506200 sw
rect 0 503200 786400 504400
rect 0 3000 3000 503200
tri 3000 503000 3200 503200 nw
tri 783200 503000 783400 503200 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 503200
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< glass >>
tri 600 503800 2400 505600 se
rect 2400 503800 784000 505600
tri 784000 503800 785800 505600 sw
rect 600 2400 2400 503800
tri 2400 503000 3200 503800 nw
tri 783200 503000 784000 503800 ne
tri 2400 2400 3200 3200 sw
tri 783200 2400 784000 3200 se
rect 784000 2400 785800 503800
tri 600 600 2400 2400 ne
rect 2400 600 784000 2400
tri 784000 600 785800 2400 nw
<< properties >>
string GDS_END 28412284
string GDS_FILE ../../gds/sealring.gds.gz
string GDS_START 104
<< end >>
