magic
tech gf180mcuD
magscale 1 10
timestamp 1764982896
<< metal1 >>
rect 12323 133 14900 185
rect 15065 133 15452 185
rect 12323 35 15345 87
rect 15511 35 15527 87
<< via1 >>
rect 14900 133 15065 185
rect 15345 35 15511 87
<< metal2 >>
rect 12368 0 12444 232
rect 13240 0 13316 232
rect 15068 187 15144 232
rect 14888 185 15144 187
rect 14888 133 14900 185
rect 15065 133 15144 185
rect 14888 131 15144 133
rect 15068 0 15144 131
rect 15256 89 15332 232
rect 15256 87 15523 89
rect 15256 35 15345 87
rect 15511 35 15523 87
rect 15256 33 15523 35
rect 15256 0 15332 33
<< end >>
