magic
tech gf180mcuD
magscale 1 5
timestamp 1764102312
<< metal2 >>
rect 0 99 950 100
rect 0 1 6 99
rect 944 1 950 99
rect 0 0 950 1
rect 1240 99 2265 100
rect 1240 1 1246 99
rect 2259 1 2265 99
rect 1240 0 2265 1
rect 2425 99 3450 100
rect 2425 1 2431 99
rect 3444 1 3450 99
rect 2425 0 3450 1
rect 3778 99 4803 100
rect 3778 1 3784 99
rect 4797 1 4803 99
rect 3778 0 4803 1
rect 4963 99 5988 100
rect 4963 1 4969 99
rect 5982 1 5988 99
rect 4963 0 5988 1
rect 6278 99 7228 100
rect 6278 1 6284 99
rect 7222 1 7228 99
rect 6278 0 7228 1
<< via2 >>
rect 6 1 944 99
rect 1246 1 2259 99
rect 2431 1 3444 99
rect 3784 1 4797 99
rect 4969 1 5982 99
rect 6284 1 7222 99
<< metal3 >>
rect 0 99 7228 100
rect 0 1 6 99
rect 944 1 1246 99
rect 2259 1 2431 99
rect 3444 1 3784 99
rect 4797 1 4969 99
rect 5982 1 6284 99
rect 7222 1 7228 99
rect 0 0 7228 1
<< via3 >>
rect 6 1 944 99
rect 1246 1 2259 99
rect 2431 1 3444 99
rect 3784 1 4797 99
rect 4969 1 5982 99
rect 6284 1 7222 99
<< metal4 >>
rect 0 99 950 100
rect 0 1 6 99
rect 944 1 950 99
rect 0 0 950 1
rect 1240 99 2265 100
rect 1240 1 1246 99
rect 2259 1 2265 99
rect 1240 0 2265 1
rect 2425 99 3450 100
rect 2425 1 2431 99
rect 3444 1 3450 99
rect 2425 0 3450 1
rect 3778 99 4803 100
rect 3778 1 3784 99
rect 4797 1 4803 99
rect 3778 0 4803 1
rect 4963 99 5988 100
rect 4963 1 4969 99
rect 5982 1 5988 99
rect 4963 0 5988 1
rect 6278 99 7228 100
rect 6278 1 6284 99
rect 7222 1 7228 99
rect 6278 0 7228 1
<< properties >>
string flatten true
<< end >>
