magic
tech gf180mcuD
magscale 1 10
timestamp 1765074735
<< checkpaint >>
rect 710929 147580 711109 160994
<< via3 >>
rect 711049 160934 711109 160994
rect 711049 160788 711109 160848
rect 711049 160641 711109 160701
rect 710929 149184 710989 149244
rect 711049 148973 711109 149033
rect 711049 148472 711109 148532
rect 711049 148330 711109 148390
rect 711049 148101 711109 148161
rect 711049 147580 711109 147640
<< end >>
