magic
tech gf180mcuD
magscale 1 10
timestamp 1765487709
<< metal2 >>
rect 89672 430768 89748 431068
rect 90193 430768 90269 431068
rect 90422 430768 90498 431068
rect 90564 430768 90640 431068
rect 90706 430768 90782 431068
rect 91066 430768 91142 431068
rect 91277 430768 91353 431068
rect 102734 430768 102810 431068
rect 102880 430768 102956 431068
rect 103026 430768 103102 431068
rect 103172 430768 103248 431068
rect 104558 430768 104634 431068
rect 104746 430768 104822 431068
rect 115472 430768 115548 431068
rect 115993 430768 116069 431068
rect 116222 430768 116298 431068
rect 116364 430768 116440 431068
rect 116506 430768 116582 431068
rect 116866 430768 116942 431068
rect 117077 430768 117153 431068
rect 128534 430768 128610 431068
rect 128680 430768 128756 431068
rect 128826 430768 128902 431068
rect 128972 430768 129048 431068
rect 130358 430768 130434 431068
rect 130546 430768 130622 431068
rect 141272 430768 141348 431068
rect 141793 430768 141869 431068
rect 142022 430768 142098 431068
rect 142164 430768 142240 431068
rect 142306 430768 142382 431068
rect 142666 430768 142742 431068
rect 142877 430768 142953 431068
rect 154334 430768 154410 431068
rect 154480 430768 154556 431068
rect 154626 430768 154702 431068
rect 154772 430768 154848 431068
rect 156158 430768 156234 431068
rect 156346 430768 156422 431068
rect 167072 430768 167148 431068
rect 167593 430768 167669 431068
rect 167822 430768 167898 431068
rect 167964 430768 168040 431068
rect 168106 430768 168182 431068
rect 168466 430768 168542 431068
rect 168677 430768 168753 431068
rect 180134 430768 180210 431068
rect 180280 430768 180356 431068
rect 180426 430768 180502 431068
rect 180572 430768 180648 431068
rect 181958 430768 182034 431068
rect 182146 430768 182222 431068
rect 244472 430768 244548 431068
rect 244993 430768 245069 431068
rect 245222 430768 245298 431068
rect 245364 430768 245440 431068
rect 245506 430768 245582 431068
rect 245866 430768 245942 431068
rect 246077 430768 246153 431068
rect 257534 430768 257610 431068
rect 257680 430768 257756 431068
rect 257826 430768 257902 431068
rect 257972 430768 258048 431068
rect 259358 430768 259434 431068
rect 259546 430768 259622 431068
rect 270272 430768 270348 431068
rect 270793 430768 270869 431068
rect 271022 430768 271098 431068
rect 271164 430768 271240 431068
rect 271306 430768 271382 431068
rect 271666 430768 271742 431068
rect 271877 430768 271953 431068
rect 283334 430768 283410 431068
rect 283480 430768 283556 431068
rect 283626 430768 283702 431068
rect 283772 430768 283848 431068
rect 285158 430768 285234 431068
rect 285346 430768 285422 431068
rect 296072 430768 296148 431068
rect 296593 430768 296669 431068
rect 296822 430768 296898 431068
rect 296964 430768 297040 431068
rect 297106 430768 297182 431068
rect 297466 430768 297542 431068
rect 297677 430768 297753 431068
rect 309134 430768 309210 431068
rect 309280 430768 309356 431068
rect 309426 430768 309502 431068
rect 309572 430768 309648 431068
rect 310958 430768 311034 431068
rect 311146 430768 311222 431068
rect 321872 430768 321948 431068
rect 322393 430768 322469 431068
rect 322622 430768 322698 431068
rect 322764 430768 322840 431068
rect 322906 430768 322982 431068
rect 323266 430768 323342 431068
rect 323477 430768 323553 431068
rect 334934 430768 335010 431068
rect 335080 430768 335156 431068
rect 335226 430768 335302 431068
rect 335372 430768 335448 431068
rect 336758 430768 336834 431068
rect 336946 430768 337022 431068
rect 347672 430768 347748 431068
rect 348193 430768 348269 431068
rect 348422 430768 348498 431068
rect 348564 430768 348640 431068
rect 348706 430768 348782 431068
rect 349066 430768 349142 431068
rect 349277 430768 349353 431068
rect 360734 430768 360810 431068
rect 360880 430768 360956 431068
rect 361026 430768 361102 431068
rect 361172 430768 361248 431068
rect 362558 430768 362634 431068
rect 362746 430768 362822 431068
rect 373472 430768 373548 431068
rect 373993 430768 374069 431068
rect 374222 430768 374298 431068
rect 374364 430768 374440 431068
rect 374506 430768 374582 431068
rect 374866 430768 374942 431068
rect 375077 430768 375153 431068
rect 386534 430768 386610 431068
rect 386680 430768 386756 431068
rect 386826 430768 386902 431068
rect 386972 430768 387048 431068
rect 388358 430768 388434 431068
rect 388546 430768 388622 431068
rect 399272 430768 399348 431068
rect 399793 430768 399869 431068
rect 400022 430768 400098 431068
rect 400164 430768 400240 431068
rect 400306 430768 400382 431068
rect 400666 430768 400742 431068
rect 400877 430768 400953 431068
rect 412334 430768 412410 431068
rect 412480 430768 412556 431068
rect 412626 430768 412702 431068
rect 412772 430768 412848 431068
rect 414158 430768 414234 431068
rect 414346 430768 414422 431068
rect 425072 430768 425148 431068
rect 425593 430768 425669 431068
rect 425822 430768 425898 431068
rect 425964 430768 426040 431068
rect 426106 430768 426182 431068
rect 426466 430768 426542 431068
rect 426677 430768 426753 431068
rect 438134 430768 438210 431068
rect 438280 430768 438356 431068
rect 438426 430768 438502 431068
rect 438572 430768 438648 431068
rect 439958 430768 440034 431068
rect 440146 430768 440222 431068
rect 450872 430768 450948 431068
rect 451393 430768 451469 431068
rect 451622 430768 451698 431068
rect 451764 430768 451840 431068
rect 451906 430768 451982 431068
rect 452266 430768 452342 431068
rect 452477 430768 452553 431068
rect 463934 430768 464010 431068
rect 464080 430768 464156 431068
rect 464226 430768 464302 431068
rect 464372 430768 464448 431068
rect 465758 430768 465834 431068
rect 465946 430768 466022 431068
rect 476672 430768 476748 431068
rect 477193 430768 477269 431068
rect 477422 430768 477498 431068
rect 477564 430768 477640 431068
rect 477706 430768 477782 431068
rect 478066 430768 478142 431068
rect 478277 430768 478353 431068
rect 489734 430768 489810 431068
rect 489880 430768 489956 431068
rect 490026 430768 490102 431068
rect 490172 430768 490248 431068
rect 491558 430768 491634 431068
rect 491746 430768 491822 431068
rect 502472 430768 502548 431068
rect 502993 430768 503069 431068
rect 503222 430768 503298 431068
rect 503364 430768 503440 431068
rect 503506 430768 503582 431068
rect 503866 430768 503942 431068
rect 504077 430768 504153 431068
rect 515534 430768 515610 431068
rect 515680 430768 515756 431068
rect 515826 430768 515902 431068
rect 515972 430768 516048 431068
rect 517358 430768 517434 431068
rect 517546 430768 517622 431068
rect 528272 430768 528348 431068
rect 528793 430768 528869 431068
rect 529022 430768 529098 431068
rect 529164 430768 529240 431068
rect 529306 430768 529382 431068
rect 529666 430768 529742 431068
rect 529877 430768 529953 431068
rect 541334 430768 541410 431068
rect 541480 430768 541556 431068
rect 541626 430768 541702 431068
rect 541772 430768 541848 431068
rect 543158 430768 543234 431068
rect 543346 430768 543422 431068
rect 605672 430768 605748 431068
rect 606193 430768 606269 431068
rect 606422 430768 606498 431068
rect 606564 430768 606640 431068
rect 606706 430768 606782 431068
rect 607066 430768 607142 431068
rect 607277 430768 607353 431068
rect 618734 430768 618810 431068
rect 618880 430768 618956 431068
rect 619026 430768 619102 431068
rect 619172 430768 619248 431068
rect 620558 430768 620634 431068
rect 620746 430768 620822 431068
rect 631472 430768 631548 431068
rect 631993 430768 632069 431068
rect 632222 430768 632298 431068
rect 632364 430768 632440 431068
rect 632506 430768 632582 431068
rect 632866 430768 632942 431068
rect 633077 430768 633153 431068
rect 644534 430768 644610 431068
rect 644680 430768 644756 431068
rect 644826 430768 644902 431068
rect 644972 430768 645048 431068
rect 646358 430768 646434 431068
rect 646546 430768 646622 431068
rect 657272 430768 657348 431068
rect 657793 430768 657869 431068
rect 658022 430768 658098 431068
rect 658164 430768 658240 431068
rect 658306 430768 658382 431068
rect 658666 430768 658742 431068
rect 658877 430768 658953 431068
rect 670334 430768 670410 431068
rect 670480 430768 670556 431068
rect 670626 430768 670702 431068
rect 670772 430768 670848 431068
rect 672158 430768 672234 431068
rect 672346 430768 672422 431068
rect 683072 430768 683148 431068
rect 683593 430768 683669 431068
rect 683822 430768 683898 431068
rect 683964 430768 684040 431068
rect 684106 430768 684182 431068
rect 684466 430768 684542 431068
rect 684677 430768 684753 431068
rect 696134 430768 696210 431068
rect 696280 430768 696356 431068
rect 696426 430768 696502 431068
rect 696572 430768 696648 431068
rect 697958 430768 698034 431068
rect 698146 430768 698222 431068
rect 74951 355724 75251 356232
rect 74951 354588 75251 355096
rect 74951 353452 75251 353960
rect 74951 352316 75251 352824
rect 74951 350776 75251 351284
rect 74951 349640 75251 350148
rect 74951 348504 75251 349012
rect 74951 347368 75251 347876
rect 74951 327524 75251 328032
rect 74951 326388 75251 326896
rect 74951 325252 75251 325760
rect 74951 324116 75251 324624
rect 74951 322576 75251 323084
rect 74951 321440 75251 321948
rect 74951 320304 75251 320812
rect 74951 319168 75251 319676
rect 74951 299324 75251 299832
rect 74951 298188 75251 298696
rect 74951 297052 75251 297560
rect 74951 295916 75251 296424
rect 74951 294376 75251 294884
rect 74951 293240 75251 293748
rect 74951 292104 75251 292612
rect 74951 290968 75251 291476
rect 74951 271124 75251 271632
rect 74951 269988 75251 270496
rect 74951 268852 75251 269360
rect 74951 267716 75251 268224
rect 74951 266176 75251 266684
rect 74951 265040 75251 265548
rect 74951 263904 75251 264412
rect 74951 262768 75251 263276
rect 89752 75102 89826 75402
rect 101858 75102 101934 75402
rect 102730 75102 102806 75402
rect 104558 75102 104634 75402
rect 104746 75102 104822 75402
rect 115552 75102 115626 75402
rect 127658 75102 127734 75402
rect 128530 75102 128606 75402
rect 130358 75102 130434 75402
rect 130546 75102 130622 75402
rect 141272 75132 141348 75432
rect 141793 75132 141869 75432
rect 142022 75132 142098 75432
rect 142164 75132 142240 75432
rect 142306 75132 142382 75432
rect 142666 75132 142742 75432
rect 142877 75132 142953 75432
rect 154334 75132 154410 75432
rect 154480 75132 154556 75432
rect 154626 75132 154702 75432
rect 154772 75132 154848 75432
rect 156158 75132 156234 75432
rect 156346 75132 156422 75432
rect 167072 75132 167148 75432
rect 167593 75132 167669 75432
rect 167822 75132 167898 75432
rect 167964 75132 168040 75432
rect 168106 75132 168182 75432
rect 168466 75132 168542 75432
rect 168677 75132 168753 75432
rect 180134 75132 180210 75432
rect 180280 75132 180356 75432
rect 180426 75132 180502 75432
rect 180572 75132 180648 75432
rect 181958 75132 182034 75432
rect 182146 75132 182222 75432
rect 244472 75132 244548 75432
rect 244993 75132 245069 75432
rect 245222 75132 245298 75432
rect 245364 75132 245440 75432
rect 245506 75132 245582 75432
rect 245866 75132 245942 75432
rect 246077 75132 246153 75432
rect 257534 75132 257610 75432
rect 257680 75132 257756 75432
rect 257826 75132 257902 75432
rect 257972 75132 258048 75432
rect 259358 75132 259434 75432
rect 259546 75132 259622 75432
rect 270272 75132 270348 75432
rect 270793 75132 270869 75432
rect 271022 75132 271098 75432
rect 271164 75132 271240 75432
rect 271306 75132 271382 75432
rect 271666 75132 271742 75432
rect 271877 75132 271953 75432
rect 283334 75132 283410 75432
rect 283480 75132 283556 75432
rect 283626 75132 283702 75432
rect 283772 75132 283848 75432
rect 285158 75132 285234 75432
rect 285346 75132 285422 75432
rect 296072 75132 296148 75432
rect 296593 75132 296669 75432
rect 296822 75132 296898 75432
rect 296964 75132 297040 75432
rect 297106 75132 297182 75432
rect 297466 75132 297542 75432
rect 297677 75132 297753 75432
rect 309134 75132 309210 75432
rect 309280 75132 309356 75432
rect 309426 75132 309502 75432
rect 309572 75132 309648 75432
rect 310958 75132 311034 75432
rect 311146 75132 311222 75432
rect 321872 75132 321948 75432
rect 322393 75132 322469 75432
rect 322622 75132 322698 75432
rect 322764 75132 322840 75432
rect 322906 75132 322982 75432
rect 323266 75132 323342 75432
rect 323477 75132 323553 75432
rect 334934 75132 335010 75432
rect 335080 75132 335156 75432
rect 335226 75132 335302 75432
rect 335372 75132 335448 75432
rect 336758 75132 336834 75432
rect 336946 75132 337022 75432
rect 347672 75132 347748 75432
rect 348193 75132 348269 75432
rect 348422 75132 348498 75432
rect 348564 75132 348640 75432
rect 348706 75132 348782 75432
rect 349066 75132 349142 75432
rect 349277 75132 349353 75432
rect 360734 75132 360810 75432
rect 360880 75132 360956 75432
rect 361026 75132 361102 75432
rect 361172 75132 361248 75432
rect 362558 75132 362634 75432
rect 362746 75132 362822 75432
rect 373472 75132 373548 75432
rect 373993 75132 374069 75432
rect 374222 75132 374298 75432
rect 374364 75132 374440 75432
rect 374506 75132 374582 75432
rect 374866 75132 374942 75432
rect 375077 75132 375153 75432
rect 386534 75132 386610 75432
rect 386680 75132 386756 75432
rect 386826 75132 386902 75432
rect 386972 75132 387048 75432
rect 388358 75132 388434 75432
rect 388546 75132 388622 75432
rect 399272 75132 399348 75432
rect 399793 75132 399869 75432
rect 400022 75132 400098 75432
rect 400164 75132 400240 75432
rect 400306 75132 400382 75432
rect 400666 75132 400742 75432
rect 400877 75132 400953 75432
rect 412334 75132 412410 75432
rect 412480 75132 412556 75432
rect 412626 75132 412702 75432
rect 412772 75132 412848 75432
rect 414158 75132 414234 75432
rect 414346 75132 414422 75432
rect 425072 75132 425148 75432
rect 425593 75132 425669 75432
rect 425822 75132 425898 75432
rect 425964 75132 426040 75432
rect 426106 75132 426182 75432
rect 426466 75132 426542 75432
rect 426677 75132 426753 75432
rect 438134 75132 438210 75432
rect 438280 75132 438356 75432
rect 438426 75132 438502 75432
rect 438572 75132 438648 75432
rect 439958 75132 440034 75432
rect 440146 75132 440222 75432
rect 450872 75132 450948 75432
rect 451393 75132 451469 75432
rect 451622 75132 451698 75432
rect 451764 75132 451840 75432
rect 451906 75132 451982 75432
rect 452266 75132 452342 75432
rect 452477 75132 452553 75432
rect 463934 75132 464010 75432
rect 464080 75132 464156 75432
rect 464226 75132 464302 75432
rect 464372 75132 464448 75432
rect 465758 75132 465834 75432
rect 465946 75132 466022 75432
rect 476672 75132 476748 75432
rect 477193 75132 477269 75432
rect 477422 75132 477498 75432
rect 477564 75132 477640 75432
rect 477706 75132 477782 75432
rect 478066 75132 478142 75432
rect 478277 75132 478353 75432
rect 489734 75132 489810 75432
rect 489880 75132 489956 75432
rect 490026 75132 490102 75432
rect 490172 75132 490248 75432
rect 491558 75132 491634 75432
rect 491746 75132 491822 75432
rect 502472 75132 502548 75432
rect 502993 75132 503069 75432
rect 503222 75132 503298 75432
rect 503364 75132 503440 75432
rect 503506 75132 503582 75432
rect 503866 75132 503942 75432
rect 504077 75132 504153 75432
rect 515534 75132 515610 75432
rect 515680 75132 515756 75432
rect 515826 75132 515902 75432
rect 515972 75132 516048 75432
rect 517358 75132 517434 75432
rect 517546 75132 517622 75432
rect 528272 75132 528348 75432
rect 528793 75132 528869 75432
rect 529022 75132 529098 75432
rect 529164 75132 529240 75432
rect 529306 75132 529382 75432
rect 529666 75132 529742 75432
rect 529877 75132 529953 75432
rect 541334 75132 541410 75432
rect 541480 75132 541556 75432
rect 541626 75132 541702 75432
rect 541772 75132 541848 75432
rect 543158 75132 543234 75432
rect 543346 75132 543422 75432
rect 605672 75132 605748 75432
rect 606193 75132 606269 75432
rect 606422 75132 606498 75432
rect 606564 75132 606640 75432
rect 606706 75132 606782 75432
rect 607066 75132 607142 75432
rect 607277 75132 607353 75432
rect 618734 75132 618810 75432
rect 618880 75132 618956 75432
rect 619026 75132 619102 75432
rect 619172 75132 619248 75432
rect 620558 75132 620634 75432
rect 620746 75132 620822 75432
rect 631472 75132 631548 75432
rect 631993 75132 632069 75432
rect 632222 75132 632298 75432
rect 632364 75132 632440 75432
rect 632506 75132 632582 75432
rect 632866 75132 632942 75432
rect 633077 75132 633153 75432
rect 644534 75132 644610 75432
rect 644680 75132 644756 75432
rect 644826 75132 644902 75432
rect 644972 75132 645048 75432
rect 646358 75132 646434 75432
rect 646546 75132 646622 75432
rect 657272 75132 657348 75432
rect 657793 75132 657869 75432
rect 658022 75132 658098 75432
rect 658164 75132 658240 75432
rect 658306 75132 658382 75432
rect 658666 75132 658742 75432
rect 658877 75132 658953 75432
rect 670334 75132 670410 75432
rect 670480 75132 670556 75432
rect 670626 75132 670702 75432
rect 670772 75132 670848 75432
rect 672158 75132 672234 75432
rect 672346 75132 672422 75432
rect 683072 75132 683148 75432
rect 683593 75132 683669 75432
rect 683822 75132 683898 75432
rect 683964 75132 684040 75432
rect 684106 75132 684182 75432
rect 684466 75132 684542 75432
rect 684677 75132 684753 75432
rect 696134 75132 696210 75432
rect 696280 75132 696356 75432
rect 696426 75132 696502 75432
rect 696572 75132 696648 75432
rect 697958 75132 698034 75432
rect 698146 75132 698222 75432
<< metal3 >>
rect 710897 360046 711197 360122
rect 710897 359858 711197 359934
rect 710897 358472 711197 358548
rect 710897 358326 711197 358402
rect 710897 358180 711197 358256
rect 710897 358034 711197 358110
rect 710897 346577 711197 346653
rect 710897 346366 711197 346442
rect 710897 346006 711197 346082
rect 710897 345864 711197 345940
rect 710897 345722 711197 345798
rect 710897 345493 711197 345569
rect 710897 344972 711197 345048
rect 710897 331846 711197 331922
rect 710897 331658 711197 331734
rect 710897 330272 711197 330348
rect 710897 330126 711197 330202
rect 710897 329980 711197 330056
rect 710897 329834 711197 329910
rect 710897 318377 711197 318453
rect 710897 318166 711197 318242
rect 710897 317806 711197 317882
rect 710897 317664 711197 317740
rect 710897 317522 711197 317598
rect 710897 317293 711197 317369
rect 710897 316772 711197 316848
rect 710897 303646 711197 303722
rect 710897 303458 711197 303534
rect 710897 302072 711197 302148
rect 710897 301926 711197 302002
rect 710897 301780 711197 301856
rect 710897 301634 711197 301710
rect 710897 290177 711197 290253
rect 710897 289966 711197 290042
rect 710897 289606 711197 289682
rect 710897 289464 711197 289540
rect 710897 289322 711197 289398
rect 710897 289093 711197 289169
rect 710897 288572 711197 288648
rect 710897 275446 711197 275522
rect 710897 275258 711197 275334
rect 710897 273872 711197 273948
rect 710897 273726 711197 273802
rect 710897 273580 711197 273656
rect 710897 273434 711197 273510
rect 710897 261977 711197 262053
rect 710897 261766 711197 261842
rect 710897 261406 711197 261482
rect 710897 261264 711197 261340
rect 710897 261122 711197 261198
rect 710897 260893 711197 260969
rect 710897 260372 711197 260448
rect 75203 247246 75503 247322
rect 710897 247246 711197 247322
rect 75203 247058 75503 247134
rect 710897 247058 711197 247134
rect 710897 245672 711197 245748
rect 710897 245526 711197 245602
rect 710897 245380 711197 245456
rect 75203 245231 75503 245307
rect 710897 245234 711197 245310
rect 75203 244358 75503 244434
rect 710897 233777 711197 233853
rect 710897 233566 711197 233642
rect 710897 233206 711197 233282
rect 710897 233064 711197 233140
rect 710897 232922 711197 232998
rect 710897 232693 711197 232769
rect 75202 232252 75503 232328
rect 710897 232172 711197 232248
rect 75203 219046 75503 219122
rect 710897 219046 711197 219122
rect 75203 218858 75503 218934
rect 710897 218858 711197 218934
rect 710897 217472 711197 217548
rect 710897 217326 711197 217402
rect 710897 217180 711197 217256
rect 75203 217031 75503 217107
rect 710897 217034 711197 217110
rect 75203 216158 75503 216234
rect 710897 205577 711197 205653
rect 710897 205366 711197 205442
rect 710897 205006 711197 205082
rect 710897 204864 711197 204940
rect 710897 204722 711197 204798
rect 710897 204493 711197 204569
rect 75203 204052 75503 204128
rect 710897 203972 711197 204048
rect 75203 190846 75503 190922
rect 710897 190846 711197 190922
rect 75203 190658 75503 190734
rect 710897 190658 711197 190734
rect 710897 189272 711197 189348
rect 710897 189126 711197 189202
rect 710897 188980 711197 189056
rect 75203 188831 75503 188907
rect 710897 188834 711197 188910
rect 75203 187958 75503 188034
rect 710897 177377 711197 177453
rect 710897 177166 711197 177242
rect 710897 176806 711197 176882
rect 710897 176664 711197 176740
rect 710897 176522 711197 176598
rect 710897 176293 711197 176369
rect 75203 175852 75503 175928
rect 710897 175772 711197 175848
rect 75203 162646 75503 162722
rect 710897 162646 711197 162722
rect 75203 162458 75503 162534
rect 710897 162458 711197 162534
rect 710897 161072 711197 161148
rect 710897 160926 711197 161002
rect 710897 160780 711197 160856
rect 75203 160631 75503 160707
rect 710897 160634 711197 160710
rect 75203 159758 75503 159834
rect 710897 149177 711197 149253
rect 710897 148966 711197 149042
rect 710897 148606 711197 148682
rect 710897 148464 711197 148540
rect 710897 148322 711197 148398
rect 710897 148093 711197 148169
rect 75203 147652 75503 147728
rect 710897 147572 711197 147648
<< metal4 >>
rect 192474 430800 194370 431000
rect 194954 430800 197000 431000
rect 197324 430800 199370 431000
rect 200030 430800 202076 431000
rect 202400 430800 204446 431000
rect 205030 430800 206926 431000
rect 218274 430800 220170 431000
rect 220754 430800 222800 431000
rect 223124 430800 225170 431000
rect 225830 430800 227876 431000
rect 228200 430800 230246 431000
rect 230830 430800 232726 431000
rect 553674 430800 555570 431000
rect 556154 430800 558200 431000
rect 558524 430800 560570 431000
rect 561230 430800 563276 431000
rect 563600 430800 565646 431000
rect 566230 430800 568126 431000
rect 579474 430800 581370 431000
rect 581954 430800 584000 431000
rect 584324 430800 586370 431000
rect 587030 430800 589076 431000
rect 589400 430800 591446 431000
rect 592030 430800 593926 431000
rect 192474 75200 194370 75400
rect 194954 75200 197000 75400
rect 197324 75200 199370 75400
rect 200030 75200 202076 75400
rect 202400 75200 204446 75400
rect 205030 75200 206926 75400
rect 218274 75200 220170 75400
rect 220754 75200 222800 75400
rect 223124 75200 225170 75400
rect 225830 75200 227876 75400
rect 228200 75200 230246 75400
rect 230830 75200 232726 75400
rect 553674 75200 555570 75400
rect 556154 75200 558200 75400
rect 558524 75200 560570 75400
rect 561230 75200 563276 75400
rect 563600 75200 565646 75400
rect 566230 75200 568126 75400
rect 579474 75200 581370 75400
rect 581954 75200 584000 75400
rect 584324 75200 586370 75400
rect 587030 75200 589076 75400
rect 589400 75200 591446 75400
rect 592030 75200 593926 75400
<< metal5 >>
rect 94032 491968 99032 496968
rect 119832 491968 124832 496968
rect 145632 491968 150632 496968
rect 171432 491968 176432 496968
rect 197232 491968 202232 496968
rect 223032 491968 228032 496968
rect 248832 491968 253832 496968
rect 274632 491968 279632 496968
rect 300432 491968 305432 496968
rect 326232 491968 331232 496968
rect 352032 491968 357032 496968
rect 377832 491968 382832 496968
rect 403632 491968 408632 496968
rect 429432 491968 434432 496968
rect 455232 491968 460232 496968
rect 481032 491968 486032 496968
rect 506832 491968 511832 496968
rect 532632 491968 537632 496968
rect 558432 491968 563432 496968
rect 584232 491968 589232 496968
rect 610032 491968 615032 496968
rect 635832 491968 640832 496968
rect 661632 491968 666632 496968
rect 687432 491968 692432 496968
rect 75200 413530 75470 415426
rect 710930 413530 711200 415426
rect 75200 410900 75470 412946
rect 710930 410900 711200 412946
rect 9200 405732 14200 410732
rect 75200 408530 75470 410576
rect 710930 408530 711200 410576
rect 75200 405824 75470 407870
rect 710930 405824 711200 407870
rect 772168 405732 777168 410732
rect 75200 403454 75470 405500
rect 710930 403454 711200 405500
rect 75200 400974 75470 402870
rect 710930 400974 711200 402870
rect 75200 385330 75470 387226
rect 710930 385330 711200 387226
rect 75200 382700 75470 384746
rect 710930 382700 711200 384746
rect 9200 377532 14200 382532
rect 75200 380330 75470 382376
rect 710930 380330 711200 382376
rect 75200 377624 75470 379670
rect 710930 377624 711200 379670
rect 772168 377532 777168 382532
rect 75200 375254 75470 377300
rect 710930 375254 711200 377300
rect 75200 372774 75470 374670
rect 710930 372774 711200 374670
rect 9200 349332 14200 354332
rect 772168 349332 777168 354332
rect 9200 321132 14200 326132
rect 772168 321132 777168 326132
rect 9200 292932 14200 297932
rect 772168 292932 777168 297932
rect 9200 264732 14200 269732
rect 772168 264732 777168 269732
rect 9200 236532 14200 241532
rect 772168 236532 777168 241532
rect 9200 208332 14200 213332
rect 772168 208332 777168 213332
rect 9200 180132 14200 185132
rect 772168 180132 777168 185132
rect 9200 151932 14200 156932
rect 772168 151932 777168 156932
rect 75200 131530 75470 133426
rect 710930 131530 711200 133426
rect 75200 128900 75470 130946
rect 710930 128900 711200 130946
rect 9200 123732 14200 128732
rect 75200 126530 75470 128576
rect 710930 126530 711200 128576
rect 75200 123824 75470 125870
rect 710930 123824 711200 125870
rect 772168 123732 777168 128732
rect 75200 121454 75470 123500
rect 710930 121454 711200 123500
rect 75200 118974 75470 120870
rect 710930 118974 711200 120870
rect 75200 103330 75470 105226
rect 710930 103330 711200 105226
rect 75200 100700 75470 102746
rect 710930 100700 711200 102746
rect 9200 95532 14200 100532
rect 75200 98330 75470 100376
rect 710930 98330 711200 100376
rect 75200 95624 75470 97670
rect 710930 95624 711200 97670
rect 772168 95532 777168 100532
rect 75200 93254 75470 95300
rect 710930 93254 711200 95300
rect 75200 90774 75470 92670
rect 710930 90774 711200 92670
rect 94032 9168 99032 14168
rect 119832 9168 124832 14168
rect 145632 9168 150632 14168
rect 171432 9168 176432 14168
rect 197232 9168 202232 14168
rect 223032 9168 228032 14168
rect 248832 9168 253832 14168
rect 274632 9168 279632 14168
rect 300432 9168 305432 14168
rect 326232 9168 331232 14168
rect 352032 9168 357032 14168
rect 377832 9168 382832 14168
rect 403632 9168 408632 14168
rect 429432 9168 434432 14168
rect 455232 9168 460232 14168
rect 481032 9168 486032 14168
rect 506832 9168 511832 14168
rect 532632 9168 537632 14168
rect 558432 9168 563432 14168
rect 584232 9168 589232 14168
rect 610032 9168 615032 14168
rect 635832 9168 640832 14168
rect 661632 9168 666632 14168
rect 687432 9168 692432 14168
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 1 5200 -1 0 274700
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_1
timestamp 1765232829
transform 0 1 5200 -1 0 302900
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_2
timestamp 1765232829
transform 0 1 5200 -1 0 359300
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_3
timestamp 1765232829
transform 0 1 5200 -1 0 331100
box -32 0 15032 70000
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 1 0 682400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_1
timestamp 1765232829
transform 1 0 656600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_2
timestamp 1765232829
transform 1 0 630800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_3
timestamp 1765232829
transform 1 0 605000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_4
timestamp 1765232829
transform 1 0 450200 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_5
timestamp 1765232829
transform 1 0 398600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_6
timestamp 1765232829
transform 1 0 476000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_7
timestamp 1765232829
transform 1 0 527600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_8
timestamp 1765232829
transform 1 0 501800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_9
timestamp 1765232829
transform 1 0 424400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_10
timestamp 1765232829
transform 0 -1 781200 1 0 175100
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_11
timestamp 1765232829
transform 0 -1 781200 1 0 146900
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_12
timestamp 1765232829
transform 0 -1 781200 1 0 203300
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_13
timestamp 1765232829
transform 0 -1 781200 1 0 231500
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_14
timestamp 1765232829
transform 1 0 269600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_15
timestamp 1765232829
transform 1 0 347000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_16
timestamp 1765232829
transform 1 0 372800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_17
timestamp 1765232829
transform 1 0 295400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_18
timestamp 1765232829
transform 1 0 321200 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_19
timestamp 1765232829
transform 1 0 243800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_20
timestamp 1765232829
transform 1 0 140600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_21
timestamp 1765232829
transform 1 0 166400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_22
timestamp 1765232829
transform 1 0 89000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_23
timestamp 1765232829
transform 1 0 140600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_24
timestamp 1765232829
transform 1 0 166400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_25
timestamp 1765232829
transform 1 0 114800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_26
timestamp 1765232829
transform 1 0 372800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_27
timestamp 1765232829
transform 1 0 295400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_28
timestamp 1765232829
transform 1 0 347000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_29
timestamp 1765232829
transform 1 0 243800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_30
timestamp 1765232829
transform 1 0 269600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_31
timestamp 1765232829
transform 1 0 321200 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_32
timestamp 1765232829
transform 0 -1 781200 1 0 287900
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_33
timestamp 1765232829
transform 0 -1 781200 1 0 259700
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_34
timestamp 1765232829
transform 0 -1 781200 1 0 316100
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_35
timestamp 1765232829
transform 0 -1 781200 1 0 344300
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_36
timestamp 1765232829
transform 1 0 501800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_37
timestamp 1765232829
transform 1 0 476000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_38
timestamp 1765232829
transform 1 0 424400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_39
timestamp 1765232829
transform 1 0 450200 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_40
timestamp 1765232829
transform 1 0 398600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_41
timestamp 1765232829
transform 1 0 527600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_42
timestamp 1765232829
transform 1 0 630800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_43
timestamp 1765232829
transform 1 0 656600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_44
timestamp 1765232829
transform 1 0 682400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_45
timestamp 1765232829
transform 1 0 605000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform -1 0 781200 0 1 5200
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_1
timestamp 1765232829
transform 1 0 5200 0 1 5200
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_2
timestamp 1765232829
transform 1 0 5200 0 -1 501000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_3
timestamp 1765232829
transform -1 0 781200 0 -1 501000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_1 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 1 0 579200 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_3
timestamp 1765232829
transform 0 1 5200 -1 0 133700
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_5
timestamp 1765232829
transform 1 0 218000 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_6
timestamp 1765232829
transform 0 -1 781200 1 0 400700
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_1 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 1 0 553400 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_2
timestamp 1765232829
transform 0 1 5200 -1 0 105500
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_5
timestamp 1765232829
transform 1 0 192200 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_7
timestamp 1765232829
transform 0 -1 781200 1 0 372500
box -32 0 15032 70000
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 118500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_1
timestamp 1765232829
transform 0 -1 781200 1 0 90200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_2
timestamp 1765232829
transform 1 0 656200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_3
timestamp 1765232829
transform 1 0 656400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_4
timestamp 1765232829
transform 1 0 681600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_5
timestamp 1765232829
transform 1 0 681800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_6
timestamp 1765232829
transform 1 0 682000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_7
timestamp 1765232829
transform 1 0 682200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_8
timestamp 1765232829
transform 1 0 709400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_9
timestamp 1765232829
transform 1 0 709600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_10
timestamp 1765232829
transform 1 0 709800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_11
timestamp 1765232829
transform 1 0 710000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_12
timestamp 1765232829
transform 1 0 656000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_13
timestamp 1765232829
transform 1 0 604200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_14
timestamp 1765232829
transform 1 0 604400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_15
timestamp 1765232829
transform 1 0 604600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_16
timestamp 1765232829
transform 1 0 604800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_17
timestamp 1765232829
transform 1 0 630000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_18
timestamp 1765232829
transform 1 0 630200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_19
timestamp 1765232829
transform 1 0 630400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_20
timestamp 1765232829
transform 1 0 630600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_21
timestamp 1765232829
transform 1 0 655800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_22
timestamp 1765232829
transform 1 0 449600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_23
timestamp 1765232829
transform 1 0 449400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_24
timestamp 1765232829
transform 1 0 424200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_25
timestamp 1765232829
transform 1 0 449800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_26
timestamp 1765232829
transform 1 0 423800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_27
timestamp 1765232829
transform 1 0 424000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_28
timestamp 1765232829
transform 1 0 450000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_29
timestamp 1765232829
transform 1 0 475200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_30
timestamp 1765232829
transform 1 0 475400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_31
timestamp 1765232829
transform 1 0 475600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_32
timestamp 1765232829
transform 1 0 475800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_33
timestamp 1765232829
transform 1 0 501000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_34
timestamp 1765232829
transform 1 0 501200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_35
timestamp 1765232829
transform 1 0 501400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_36
timestamp 1765232829
transform 1 0 501600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_37
timestamp 1765232829
transform 1 0 526800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_38
timestamp 1765232829
transform 1 0 423600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_39
timestamp 1765232829
transform 1 0 397800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_40
timestamp 1765232829
transform 1 0 398000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_41
timestamp 1765232829
transform 1 0 398200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_42
timestamp 1765232829
transform 1 0 398400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_43
timestamp 1765232829
transform 1 0 527000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_44
timestamp 1765232829
transform 1 0 527400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_45
timestamp 1765232829
transform 1 0 527200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_46
timestamp 1765232829
transform 1 0 552600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_47
timestamp 1765232829
transform 1 0 552800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_48
timestamp 1765232829
transform 1 0 553000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_49
timestamp 1765232829
transform 1 0 553200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_50
timestamp 1765232829
transform 1 0 578400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_51
timestamp 1765232829
transform 1 0 578600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_52
timestamp 1765232829
transform 1 0 578800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_53
timestamp 1765232829
transform 1 0 579000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_54
timestamp 1765232829
transform 0 -1 781200 1 0 146700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_55
timestamp 1765232829
transform 0 -1 781200 1 0 174900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_56
timestamp 1765232829
transform 0 -1 781200 1 0 203100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_57
timestamp 1765232829
transform 0 -1 781200 1 0 231300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_58
timestamp 1765232829
transform 1 0 268800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_59
timestamp 1765232829
transform 1 0 321000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_60
timestamp 1765232829
transform 1 0 320800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_61
timestamp 1765232829
transform 1 0 320600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_62
timestamp 1765232829
transform 1 0 320400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_63
timestamp 1765232829
transform 1 0 346200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_64
timestamp 1765232829
transform 1 0 346400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_65
timestamp 1765232829
transform 1 0 346600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_66
timestamp 1765232829
transform 1 0 346800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_67
timestamp 1765232829
transform 1 0 372000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_68
timestamp 1765232829
transform 1 0 269000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_69
timestamp 1765232829
transform 1 0 295200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_70
timestamp 1765232829
transform 1 0 372400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_71
timestamp 1765232829
transform 1 0 372600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_72
timestamp 1765232829
transform 1 0 295000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_73
timestamp 1765232829
transform 1 0 294800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_74
timestamp 1765232829
transform 1 0 294600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_75
timestamp 1765232829
transform 1 0 269400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_76
timestamp 1765232829
transform 1 0 269200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_77
timestamp 1765232829
transform 1 0 372200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_78
timestamp 1765232829
transform 1 0 217800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_79
timestamp 1765232829
transform 1 0 217200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_80
timestamp 1765232829
transform 1 0 217600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_81
timestamp 1765232829
transform 1 0 217400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_82
timestamp 1765232829
transform 1 0 243600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_83
timestamp 1765232829
transform 1 0 243400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_84
timestamp 1765232829
transform 1 0 243200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_85
timestamp 1765232829
transform 1 0 243000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_86
timestamp 1765232829
transform 0 1 5200 -1 0 118700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_87
timestamp 1765232829
transform 0 1 5200 -1 0 90400
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_88
timestamp 1765232829
transform 1 0 88200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_89
timestamp 1765232829
transform 1 0 88400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_90
timestamp 1765232829
transform 1 0 88600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_91
timestamp 1765232829
transform 1 0 88800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_92
timestamp 1765232829
transform 1 0 139800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_93
timestamp 1765232829
transform 1 0 140000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_94
timestamp 1765232829
transform 1 0 140400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_95
timestamp 1765232829
transform 1 0 165600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_96
timestamp 1765232829
transform 1 0 165800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_97
timestamp 1765232829
transform 1 0 166000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_98
timestamp 1765232829
transform 1 0 166200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_99
timestamp 1765232829
transform 1 0 191400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_100
timestamp 1765232829
transform 1 0 191600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_101
timestamp 1765232829
transform 1 0 191800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_102
timestamp 1765232829
transform 1 0 192000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_103
timestamp 1765232829
transform 1 0 140200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_104
timestamp 1765232829
transform 1 0 114000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_105
timestamp 1765232829
transform 1 0 114400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_106
timestamp 1765232829
transform 1 0 114600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_107
timestamp 1765232829
transform 1 0 114200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_108
timestamp 1765232829
transform 0 1 5200 -1 0 175100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_109
timestamp 1765232829
transform 0 1 5200 -1 0 146900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_110
timestamp 1765232829
transform 0 1 5200 -1 0 231500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_111
timestamp 1765232829
transform 0 1 5200 -1 0 203300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_112
timestamp 1765232829
transform 0 1 5200 -1 0 287900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_113
timestamp 1765232829
transform 0 1 5200 -1 0 259700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_114
timestamp 1765232829
transform 0 1 5200 -1 0 344300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_115
timestamp 1765232829
transform 0 1 5200 -1 0 372500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_116
timestamp 1765232829
transform 0 1 5200 -1 0 316100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_117
timestamp 1765232829
transform 0 1 5200 -1 0 429900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_118
timestamp 1765232829
transform 0 1 5200 -1 0 400700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_119
timestamp 1765232829
transform 1 0 165600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_120
timestamp 1765232829
transform 1 0 114400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_121
timestamp 1765232829
transform 1 0 88800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_122
timestamp 1765232829
transform 1 0 88600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_123
timestamp 1765232829
transform 1 0 88400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_124
timestamp 1765232829
transform 1 0 114600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_125
timestamp 1765232829
transform 1 0 88200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_126
timestamp 1765232829
transform 1 0 139800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_127
timestamp 1765232829
transform 1 0 140000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_128
timestamp 1765232829
transform 1 0 140200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_129
timestamp 1765232829
transform 1 0 140400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_130
timestamp 1765232829
transform 1 0 191400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_131
timestamp 1765232829
transform 1 0 191600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_132
timestamp 1765232829
transform 1 0 166200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_133
timestamp 1765232829
transform 1 0 191800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_134
timestamp 1765232829
transform 1 0 166000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_135
timestamp 1765232829
transform 1 0 165800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_136
timestamp 1765232829
transform 1 0 192000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_137
timestamp 1765232829
transform 1 0 114000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_138
timestamp 1765232829
transform 1 0 114200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_139
timestamp 1765232829
transform 1 0 321000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_140
timestamp 1765232829
transform 1 0 269000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_141
timestamp 1765232829
transform 1 0 320800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_142
timestamp 1765232829
transform 1 0 269400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_143
timestamp 1765232829
transform 1 0 294600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_144
timestamp 1765232829
transform 1 0 294800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_145
timestamp 1765232829
transform 1 0 295000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_146
timestamp 1765232829
transform 1 0 295200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_147
timestamp 1765232829
transform 1 0 320400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_148
timestamp 1765232829
transform 1 0 320600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_149
timestamp 1765232829
transform 1 0 269200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_150
timestamp 1765232829
transform 1 0 346200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_151
timestamp 1765232829
transform 1 0 243400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_152
timestamp 1765232829
transform 1 0 243200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_153
timestamp 1765232829
transform 1 0 243000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_154
timestamp 1765232829
transform 1 0 268800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_155
timestamp 1765232829
transform 1 0 217200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_156
timestamp 1765232829
transform 1 0 217800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_157
timestamp 1765232829
transform 1 0 217600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_158
timestamp 1765232829
transform 1 0 217400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_159
timestamp 1765232829
transform 1 0 243600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_160
timestamp 1765232829
transform 1 0 346400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_161
timestamp 1765232829
transform 1 0 372600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_162
timestamp 1765232829
transform 1 0 372400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_163
timestamp 1765232829
transform 1 0 372200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_164
timestamp 1765232829
transform 1 0 372000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_165
timestamp 1765232829
transform 1 0 346800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_166
timestamp 1765232829
transform 1 0 346600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_167
timestamp 1765232829
transform 0 -1 781200 1 0 287700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_168
timestamp 1765232829
transform 0 -1 781200 1 0 259500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_169
timestamp 1765232829
transform 0 -1 781200 1 0 315900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_170
timestamp 1765232829
transform 0 -1 781200 1 0 344100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_171
timestamp 1765232829
transform 0 -1 781200 1 0 372300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_172
timestamp 1765232829
transform 1 0 579000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_173
timestamp 1765232829
transform 1 0 450000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_174
timestamp 1765232829
transform 1 0 449800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_175
timestamp 1765232829
transform 1 0 578400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_176
timestamp 1765232829
transform 1 0 578600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_177
timestamp 1765232829
transform 1 0 527400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_178
timestamp 1765232829
transform 1 0 527200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_179
timestamp 1765232829
transform 1 0 527000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_180
timestamp 1765232829
transform 1 0 526800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_181
timestamp 1765232829
transform 1 0 552600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_182
timestamp 1765232829
transform 1 0 501600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_183
timestamp 1765232829
transform 1 0 552800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_184
timestamp 1765232829
transform 1 0 449600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_185
timestamp 1765232829
transform 1 0 501200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_186
timestamp 1765232829
transform 1 0 501000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_187
timestamp 1765232829
transform 1 0 553000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_188
timestamp 1765232829
transform 1 0 553200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_189
timestamp 1765232829
transform 1 0 578800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_190
timestamp 1765232829
transform 1 0 475800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_191
timestamp 1765232829
transform 1 0 475600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_192
timestamp 1765232829
transform 1 0 475400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_193
timestamp 1765232829
transform 1 0 475200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_194
timestamp 1765232829
transform 1 0 501400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_195
timestamp 1765232829
transform 1 0 449400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_196
timestamp 1765232829
transform 1 0 424200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_197
timestamp 1765232829
transform 1 0 424000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_198
timestamp 1765232829
transform 1 0 423800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_199
timestamp 1765232829
transform 1 0 423600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_200
timestamp 1765232829
transform 1 0 398400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_201
timestamp 1765232829
transform 1 0 398000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_202
timestamp 1765232829
transform 1 0 397800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_203
timestamp 1765232829
transform 1 0 398200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_204
timestamp 1765232829
transform 0 -1 781200 1 0 429700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_205
timestamp 1765232829
transform 0 -1 781200 1 0 400500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_206
timestamp 1765232829
transform 1 0 681600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_207
timestamp 1765232829
transform 1 0 682200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_208
timestamp 1765232829
transform 1 0 682000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_209
timestamp 1765232829
transform 1 0 630000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_210
timestamp 1765232829
transform 1 0 681800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_211
timestamp 1765232829
transform 1 0 656400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_212
timestamp 1765232829
transform 1 0 709800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_213
timestamp 1765232829
transform 1 0 656200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_214
timestamp 1765232829
transform 1 0 656000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_215
timestamp 1765232829
transform 1 0 655800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_216
timestamp 1765232829
transform 1 0 604800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_217
timestamp 1765232829
transform 1 0 604200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_218
timestamp 1765232829
transform 1 0 604400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_219
timestamp 1765232829
transform 1 0 604600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_220
timestamp 1765232829
transform 1 0 710000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_221
timestamp 1765232829
transform 1 0 630200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_222
timestamp 1765232829
transform 1 0 630400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_223
timestamp 1765232829
transform 1 0 709400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_224
timestamp 1765232829
transform 1 0 630600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_225
timestamp 1765232829
transform 1 0 709600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 117500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_1
timestamp 1765232829
transform 0 -1 781200 1 0 173900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_2
timestamp 1765232829
transform 0 -1 781200 1 0 145700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_3
timestamp 1765232829
transform 0 -1 781200 1 0 202100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_4
timestamp 1765232829
transform 0 -1 781200 1 0 230300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_5
timestamp 1765232829
transform 0 1 5200 -1 0 118500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_6
timestamp 1765232829
transform 0 1 5200 -1 0 174900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_7
timestamp 1765232829
transform 0 1 5200 -1 0 146700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_8
timestamp 1765232829
transform 0 1 5200 -1 0 203100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_9
timestamp 1765232829
transform 0 1 5200 -1 0 231300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_10
timestamp 1765232829
transform 0 1 5200 -1 0 259500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_11
timestamp 1765232829
transform 0 1 5200 -1 0 287700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_12
timestamp 1765232829
transform 0 1 5200 -1 0 372300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_13
timestamp 1765232829
transform 0 1 5200 -1 0 344100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_14
timestamp 1765232829
transform 0 1 5200 -1 0 315900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_15
timestamp 1765232829
transform 0 1 5200 -1 0 400500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_16
timestamp 1765232829
transform 0 -1 781200 1 0 258500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_17
timestamp 1765232829
transform 0 -1 781200 1 0 286700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_18
timestamp 1765232829
transform 0 -1 781200 1 0 371300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_19
timestamp 1765232829
transform 0 -1 781200 1 0 343100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_20
timestamp 1765232829
transform 0 -1 781200 1 0 314900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_21
timestamp 1765232829
transform 0 -1 781200 1 0 399500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 115500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1
timestamp 1765232829
transform 0 -1 781200 1 0 105500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_2
timestamp 1765232829
transform 0 -1 781200 1 0 82200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_3
timestamp 1765232829
transform 0 -1 781200 1 0 107500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_4
timestamp 1765232829
transform 0 -1 781200 1 0 80200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_5
timestamp 1765232829
transform 0 -1 781200 1 0 78200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_6
timestamp 1765232829
transform 0 -1 781200 1 0 86200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_7
timestamp 1765232829
transform 0 -1 781200 1 0 76200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_8
timestamp 1765232829
transform 0 -1 781200 1 0 113500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_9
timestamp 1765232829
transform 0 -1 781200 1 0 111500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_10
timestamp 1765232829
transform 0 -1 781200 1 0 88200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_11
timestamp 1765232829
transform 0 -1 781200 1 0 84200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_12
timestamp 1765232829
transform 0 -1 781200 1 0 109500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_14
timestamp 1765232829
transform 1 0 679600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_15
timestamp 1765232829
transform 1 0 677600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_16
timestamp 1765232829
transform 1 0 675600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_17
timestamp 1765232829
transform 1 0 673600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_18
timestamp 1765232829
transform 1 0 626000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_19
timestamp 1765232829
transform 1 0 624000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_20
timestamp 1765232829
transform 1 0 628000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_21
timestamp 1765232829
transform 1 0 622000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_23
timestamp 1765232829
transform 1 0 602200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_24
timestamp 1765232829
transform 1 0 600200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_26
timestamp 1765232829
transform 1 0 598200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_27
timestamp 1765232829
transform 1 0 596200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_28
timestamp 1765232829
transform 1 0 594200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_29
timestamp 1765232829
transform 1 0 647800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_30
timestamp 1765232829
transform 1 0 649800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_31
timestamp 1765232829
transform 1 0 651800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_32
timestamp 1765232829
transform 1 0 653800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_33
timestamp 1765232829
transform 1 0 703400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_34
timestamp 1765232829
transform 1 0 705400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_35
timestamp 1765232829
transform 1 0 699400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_37
timestamp 1765232829
transform 1 0 701400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_38
timestamp 1765232829
transform 1 0 707400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_39
timestamp 1765232829
transform 1 0 568400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_40
timestamp 1765232829
transform 1 0 471200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_41
timestamp 1765232829
transform 1 0 570400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_42
timestamp 1765232829
transform 1 0 497000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_43
timestamp 1765232829
transform 1 0 574400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_44
timestamp 1765232829
transform 1 0 550600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_45
timestamp 1765232829
transform 1 0 447400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_46
timestamp 1765232829
transform 1 0 495000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_48
timestamp 1765232829
transform 1 0 467200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_49
timestamp 1765232829
transform 1 0 469200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_50
timestamp 1765232829
transform 1 0 445400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_51
timestamp 1765232829
transform 1 0 576400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_52
timestamp 1765232829
transform 1 0 493000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_53
timestamp 1765232829
transform 1 0 473200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_55
timestamp 1765232829
transform 1 0 415600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_56
timestamp 1765232829
transform 1 0 417600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_57
timestamp 1765232829
transform 1 0 419600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_60
timestamp 1765232829
transform 1 0 524800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_61
timestamp 1765232829
transform 1 0 572400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_62
timestamp 1765232829
transform 1 0 395800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_63
timestamp 1765232829
transform 1 0 393800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_64
timestamp 1765232829
transform 1 0 520800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_66
timestamp 1765232829
transform 1 0 441400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_67
timestamp 1765232829
transform 1 0 548600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_68
timestamp 1765232829
transform 1 0 499000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_69
timestamp 1765232829
transform 1 0 443400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_70
timestamp 1765232829
transform 1 0 518800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_72
timestamp 1765232829
transform 1 0 546600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_73
timestamp 1765232829
transform 1 0 522800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_74
timestamp 1765232829
transform 1 0 421600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_75
timestamp 1765232829
transform 1 0 544600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_76
timestamp 1765232829
transform 0 -1 781200 1 0 165900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_77
timestamp 1765232829
transform 0 -1 781200 1 0 163900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_79
timestamp 1765232829
transform 0 -1 781200 1 0 141700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_80
timestamp 1765232829
transform 0 -1 781200 1 0 139700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_81
timestamp 1765232829
transform 0 -1 781200 1 0 137700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_82
timestamp 1765232829
transform 0 -1 781200 1 0 135700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_83
timestamp 1765232829
transform 0 -1 781200 1 0 133700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_84
timestamp 1765232829
transform 0 -1 781200 1 0 143700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_85
timestamp 1765232829
transform 0 -1 781200 1 0 169900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_86
timestamp 1765232829
transform 0 -1 781200 1 0 171900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_87
timestamp 1765232829
transform 0 -1 781200 1 0 167900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_88
timestamp 1765232829
transform 0 -1 781200 1 0 224300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_89
timestamp 1765232829
transform 0 -1 781200 1 0 226300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_90
timestamp 1765232829
transform 0 -1 781200 1 0 222300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_91
timestamp 1765232829
transform 0 -1 781200 1 0 220300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_92
timestamp 1765232829
transform 0 -1 781200 1 0 228300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_95
timestamp 1765232829
transform 0 -1 781200 1 0 248500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_96
timestamp 1765232829
transform 0 -1 781200 1 0 200100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_97
timestamp 1765232829
transform 0 -1 781200 1 0 198100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_98
timestamp 1765232829
transform 0 -1 781200 1 0 196100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_99
timestamp 1765232829
transform 0 -1 781200 1 0 194100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_100
timestamp 1765232829
transform 0 -1 781200 1 0 192100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_101
timestamp 1765232829
transform 0 -1 781200 1 0 250500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_104
timestamp 1765232829
transform 1 0 260800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_105
timestamp 1765232829
transform 1 0 237000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_107
timestamp 1765232829
transform 1 0 314400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_108
timestamp 1765232829
transform 1 0 312400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_109
timestamp 1765232829
transform 1 0 235000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_110
timestamp 1765232829
transform 1 0 286600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_111
timestamp 1765232829
transform 1 0 288600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_112
timestamp 1765232829
transform 1 0 290600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_114
timestamp 1765232829
transform 1 0 266800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_115
timestamp 1765232829
transform 1 0 241000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_116
timestamp 1765232829
transform 1 0 292600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_117
timestamp 1765232829
transform 1 0 264800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_118
timestamp 1765232829
transform 1 0 262800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_119
timestamp 1765232829
transform 1 0 239000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_120
timestamp 1765232829
transform 1 0 233000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_122
timestamp 1765232829
transform 1 0 366000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_123
timestamp 1765232829
transform 1 0 318400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_124
timestamp 1765232829
transform 1 0 389800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_125
timestamp 1765232829
transform 1 0 364000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_127
timestamp 1765232829
transform 1 0 211200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_128
timestamp 1765232829
transform 1 0 209200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_129
timestamp 1765232829
transform 1 0 344200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_130
timestamp 1765232829
transform 1 0 207200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_131
timestamp 1765232829
transform 1 0 342200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_132
timestamp 1765232829
transform 1 0 340200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_133
timestamp 1765232829
transform 1 0 213200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_134
timestamp 1765232829
transform 1 0 338200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_135
timestamp 1765232829
transform 1 0 368000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_136
timestamp 1765232829
transform 1 0 316400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_137
timestamp 1765232829
transform 1 0 370000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_139
timestamp 1765232829
transform 1 0 215200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_140
timestamp 1765232829
transform 0 1 5200 -1 0 82200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_141
timestamp 1765232829
transform 0 1 5200 -1 0 84200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_142
timestamp 1765232829
transform 0 1 5200 -1 0 80200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_143
timestamp 1765232829
transform 0 1 5200 -1 0 88200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_144
timestamp 1765232829
transform 0 1 5200 -1 0 86200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_145
timestamp 1765232829
transform 0 1 5200 -1 0 78200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_146
timestamp 1765232829
transform 0 1 5200 -1 0 90200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_147
timestamp 1765232829
transform 0 1 5200 -1 0 107500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_148
timestamp 1765232829
transform 0 1 5200 -1 0 109500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_149
timestamp 1765232829
transform 0 1 5200 -1 0 111500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_150
timestamp 1765232829
transform 0 1 5200 -1 0 113500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_151
timestamp 1765232829
transform 0 1 5200 -1 0 115500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_152
timestamp 1765232829
transform 0 1 5200 -1 0 117500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_153
timestamp 1765232829
transform 1 0 106000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_155
timestamp 1765232829
transform 1 0 108000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_156
timestamp 1765232829
transform 1 0 112000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_157
timestamp 1765232829
transform 1 0 110000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_158
timestamp 1765232829
transform 1 0 163600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_159
timestamp 1765232829
transform 1 0 161600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_160
timestamp 1765232829
transform 1 0 159600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_161
timestamp 1765232829
transform 1 0 157600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_162
timestamp 1765232829
transform 1 0 131800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_164
timestamp 1765232829
transform 1 0 86200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_165
timestamp 1765232829
transform 1 0 137800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_166
timestamp 1765232829
transform 1 0 135800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_167
timestamp 1765232829
transform 1 0 133800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_168
timestamp 1765232829
transform 1 0 187400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_169
timestamp 1765232829
transform 1 0 185400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_170
timestamp 1765232829
transform 1 0 183400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_172
timestamp 1765232829
transform 1 0 189400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_173
timestamp 1765232829
transform 1 0 78200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_174
timestamp 1765232829
transform 1 0 76200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_175
timestamp 1765232829
transform 1 0 84200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_176
timestamp 1765232829
transform 1 0 80200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_178
timestamp 1765232829
transform 1 0 82200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_179
timestamp 1765232829
transform 0 1 5200 -1 0 167900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_180
timestamp 1765232829
transform 0 1 5200 -1 0 169900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_181
timestamp 1765232829
transform 0 1 5200 -1 0 171900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_182
timestamp 1765232829
transform 0 1 5200 -1 0 173900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_183
timestamp 1765232829
transform 0 1 5200 -1 0 135700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_184
timestamp 1765232829
transform 0 1 5200 -1 0 165900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_185
timestamp 1765232829
transform 0 1 5200 -1 0 137700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_186
timestamp 1765232829
transform 0 1 5200 -1 0 139700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_187
timestamp 1765232829
transform 0 1 5200 -1 0 141700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_188
timestamp 1765232829
transform 0 1 5200 -1 0 143700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_189
timestamp 1765232829
transform 0 1 5200 -1 0 145700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_191
timestamp 1765232829
transform 0 1 5200 -1 0 194100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_192
timestamp 1765232829
transform 0 1 5200 -1 0 196100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_193
timestamp 1765232829
transform 0 1 5200 -1 0 226300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_194
timestamp 1765232829
transform 0 1 5200 -1 0 198100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_195
timestamp 1765232829
transform 0 1 5200 -1 0 200100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_196
timestamp 1765232829
transform 0 1 5200 -1 0 202100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_198
timestamp 1765232829
transform 0 1 5200 -1 0 222300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_199
timestamp 1765232829
transform 0 1 5200 -1 0 224300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_200
timestamp 1765232829
transform 0 1 5200 -1 0 250500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_201
timestamp 1765232829
transform 0 1 5200 -1 0 252500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_202
timestamp 1765232829
transform 0 1 5200 -1 0 228300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_203
timestamp 1765232829
transform 0 1 5200 -1 0 230300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_206
timestamp 1765232829
transform 0 1 5200 -1 0 284700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_207
timestamp 1765232829
transform 0 1 5200 -1 0 282700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_208
timestamp 1765232829
transform 0 1 5200 -1 0 280700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_209
timestamp 1765232829
transform 0 1 5200 -1 0 278700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_210
timestamp 1765232829
transform 0 1 5200 -1 0 276700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_211
timestamp 1765232829
transform 0 1 5200 -1 0 258500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_212
timestamp 1765232829
transform 0 1 5200 -1 0 256500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_213
timestamp 1765232829
transform 0 1 5200 -1 0 286700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_214
timestamp 1765232829
transform 0 1 5200 -1 0 314900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_215
timestamp 1765232829
transform 0 1 5200 -1 0 312900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_216
timestamp 1765232829
transform 0 1 5200 -1 0 310900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_217
timestamp 1765232829
transform 0 1 5200 -1 0 308900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_218
timestamp 1765232829
transform 0 1 5200 -1 0 306900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_219
timestamp 1765232829
transform 0 1 5200 -1 0 304900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_220
timestamp 1765232829
transform 0 1 5200 -1 0 333100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_221
timestamp 1765232829
transform 0 1 5200 -1 0 335100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_222
timestamp 1765232829
transform 0 1 5200 -1 0 371300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_223
timestamp 1765232829
transform 0 1 5200 -1 0 369300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_224
timestamp 1765232829
transform 0 1 5200 -1 0 367300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_225
timestamp 1765232829
transform 0 1 5200 -1 0 365300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_226
timestamp 1765232829
transform 0 1 5200 -1 0 363300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_227
timestamp 1765232829
transform 0 1 5200 -1 0 343100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_228
timestamp 1765232829
transform 0 1 5200 -1 0 341100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_229
timestamp 1765232829
transform 0 1 5200 -1 0 361300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_230
timestamp 1765232829
transform 0 1 5200 -1 0 339100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_231
timestamp 1765232829
transform 0 1 5200 -1 0 337100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_232
timestamp 1765232829
transform 0 1 5200 -1 0 423700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_233
timestamp 1765232829
transform 0 1 5200 -1 0 425700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_234
timestamp 1765232829
transform 0 1 5200 -1 0 427700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_235
timestamp 1765232829
transform 0 1 5200 -1 0 419700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_236
timestamp 1765232829
transform 0 1 5200 -1 0 429700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_237
timestamp 1765232829
transform 0 1 5200 -1 0 417700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_238
timestamp 1765232829
transform 0 1 5200 -1 0 399500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_239
timestamp 1765232829
transform 0 1 5200 -1 0 395500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_240
timestamp 1765232829
transform 0 1 5200 -1 0 393500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_241
timestamp 1765232829
transform 0 1 5200 -1 0 391500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_242
timestamp 1765232829
transform 0 1 5200 -1 0 389500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_243
timestamp 1765232829
transform 0 1 5200 -1 0 397500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_244
timestamp 1765232829
transform 0 1 5200 -1 0 421700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_245
timestamp 1765232829
transform 1 0 131800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_246
timestamp 1765232829
transform 1 0 133800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_248
timestamp 1765232829
transform 1 0 135800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_249
timestamp 1765232829
transform 1 0 76200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_250
timestamp 1765232829
transform 1 0 78200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_251
timestamp 1765232829
transform 1 0 80200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_252
timestamp 1765232829
transform 1 0 82200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_253
timestamp 1765232829
transform 1 0 84200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_254
timestamp 1765232829
transform 1 0 86200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_255
timestamp 1765232829
transform 1 0 189400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_256
timestamp 1765232829
transform 1 0 185400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_257
timestamp 1765232829
transform 1 0 183400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_259
timestamp 1765232829
transform 1 0 159600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_260
timestamp 1765232829
transform 1 0 163600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_261
timestamp 1765232829
transform 1 0 161600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_262
timestamp 1765232829
transform 1 0 187400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_263
timestamp 1765232829
transform 1 0 137800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_265
timestamp 1765232829
transform 1 0 157600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_267
timestamp 1765232829
transform 1 0 106000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_268
timestamp 1765232829
transform 1 0 108000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_269
timestamp 1765232829
transform 1 0 110000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_270
timestamp 1765232829
transform 1 0 112000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_272
timestamp 1765232829
transform 1 0 389800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_273
timestamp 1765232829
transform 1 0 266800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_274
timestamp 1765232829
transform 1 0 264800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_275
timestamp 1765232829
transform 1 0 262800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_276
timestamp 1765232829
transform 1 0 318400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_277
timestamp 1765232829
transform 1 0 316400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_278
timestamp 1765232829
transform 1 0 314400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_279
timestamp 1765232829
transform 1 0 312400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_281
timestamp 1765232829
transform 1 0 338200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_282
timestamp 1765232829
transform 1 0 292600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_283
timestamp 1765232829
transform 1 0 340200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_284
timestamp 1765232829
transform 1 0 290600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_285
timestamp 1765232829
transform 1 0 342200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_286
timestamp 1765232829
transform 1 0 344200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_288
timestamp 1765232829
transform 1 0 364000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_289
timestamp 1765232829
transform 1 0 366000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_290
timestamp 1765232829
transform 1 0 288600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_291
timestamp 1765232829
transform 1 0 368000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_292
timestamp 1765232829
transform 1 0 370000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_293
timestamp 1765232829
transform 1 0 286600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_295
timestamp 1765232829
transform 1 0 213200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_296
timestamp 1765232829
transform 1 0 211200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_297
timestamp 1765232829
transform 1 0 209200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_298
timestamp 1765232829
transform 1 0 207200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_299
timestamp 1765232829
transform 1 0 260800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_301
timestamp 1765232829
transform 1 0 241000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_302
timestamp 1765232829
transform 1 0 239000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_303
timestamp 1765232829
transform 1 0 237000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_304
timestamp 1765232829
transform 1 0 235000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_305
timestamp 1765232829
transform 1 0 233000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_306
timestamp 1765232829
transform 1 0 215200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_308
timestamp 1765232829
transform 0 -1 781200 1 0 282700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_309
timestamp 1765232829
transform 0 -1 781200 1 0 284700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10_310x
timestamp 1765487709
transform 0 -1 781200 1 0 302900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_311
timestamp 1765232829
transform 0 -1 781200 1 0 304900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_312
timestamp 1765232829
transform 0 -1 781200 1 0 306900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_313
timestamp 1765232829
transform 0 -1 781200 1 0 308900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_314
timestamp 1765232829
transform 0 -1 781200 1 0 310900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_315
timestamp 1765232829
transform 0 -1 781200 1 0 312900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_316
timestamp 1765232829
transform 0 -1 781200 1 0 254500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_317
timestamp 1765232829
transform 0 -1 781200 1 0 256500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_319
timestamp 1765232829
transform 0 -1 781200 1 0 276700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_320
timestamp 1765232829
transform 0 -1 781200 1 0 278700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_321
timestamp 1765232829
transform 0 -1 781200 1 0 280700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_322
timestamp 1765232829
transform 0 -1 781200 1 0 361300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_324
timestamp 1765232829
transform 0 -1 781200 1 0 333100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_325
timestamp 1765232829
transform 0 -1 781200 1 0 335100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_326
timestamp 1765232829
transform 0 -1 781200 1 0 337100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_327
timestamp 1765232829
transform 0 -1 781200 1 0 369300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_328
timestamp 1765232829
transform 0 -1 781200 1 0 367300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_329
timestamp 1765232829
transform 0 -1 781200 1 0 365300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_330
timestamp 1765232829
transform 0 -1 781200 1 0 363300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_332
timestamp 1765232829
transform 0 -1 781200 1 0 341100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_333
timestamp 1765232829
transform 0 -1 781200 1 0 339100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_334
timestamp 1765232829
transform 1 0 393800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_335
timestamp 1765232829
transform 1 0 395800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_337
timestamp 1765232829
transform 1 0 415600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_338
timestamp 1765232829
transform 1 0 417600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_339
timestamp 1765232829
transform 1 0 419600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_340
timestamp 1765232829
transform 1 0 421600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_342
timestamp 1765232829
transform 1 0 441400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_343
timestamp 1765232829
transform 1 0 443400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_344
timestamp 1765232829
transform 1 0 447400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_346
timestamp 1765232829
transform 1 0 467200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_347
timestamp 1765232829
transform 1 0 469200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_348
timestamp 1765232829
transform 1 0 471200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_349
timestamp 1765232829
transform 1 0 473200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_351
timestamp 1765232829
transform 1 0 493000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_352
timestamp 1765232829
transform 1 0 495000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_353
timestamp 1765232829
transform 1 0 497000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_354
timestamp 1765232829
transform 1 0 499000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_356
timestamp 1765232829
transform 1 0 518800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_357
timestamp 1765232829
transform 1 0 445400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_358
timestamp 1765232829
transform 1 0 520800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_359
timestamp 1765232829
transform 1 0 522800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_360
timestamp 1765232829
transform 1 0 524800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_362
timestamp 1765232829
transform 1 0 544600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_363
timestamp 1765232829
transform 1 0 546600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_364
timestamp 1765232829
transform 1 0 548600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_365
timestamp 1765232829
transform 1 0 550600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_366
timestamp 1765232829
transform 1 0 568400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_367
timestamp 1765232829
transform 1 0 570400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_368
timestamp 1765232829
transform 1 0 574400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_369
timestamp 1765232829
transform 1 0 576400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_370
timestamp 1765232829
transform 1 0 572400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_371
timestamp 1765232829
transform 0 -1 781200 1 0 389500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_372
timestamp 1765232829
transform 0 -1 781200 1 0 391500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_373
timestamp 1765232829
transform 0 -1 781200 1 0 423700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_374
timestamp 1765232829
transform 0 -1 781200 1 0 421700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_375
timestamp 1765232829
transform 0 -1 781200 1 0 387500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_376
timestamp 1765232829
transform 0 -1 781200 1 0 417700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_377
timestamp 1765232829
transform 0 -1 781200 1 0 419700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_378
timestamp 1765232829
transform 0 -1 781200 1 0 397500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_379
timestamp 1765232829
transform 0 -1 781200 1 0 415700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_380
timestamp 1765232829
transform 0 -1 781200 1 0 395500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_381
timestamp 1765232829
transform 0 -1 781200 1 0 425700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_382
timestamp 1765232829
transform 0 -1 781200 1 0 393500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_383
timestamp 1765232829
transform 0 -1 781200 1 0 427700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_384
timestamp 1765232829
transform 1 0 707400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_385
timestamp 1765232829
transform 1 0 705400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_386
timestamp 1765232829
transform 1 0 703400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_387
timestamp 1765232829
transform 1 0 602200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_388
timestamp 1765232829
transform 1 0 701400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_390
timestamp 1765232829
transform 1 0 622000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_391
timestamp 1765232829
transform 1 0 624000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_392
timestamp 1765232829
transform 1 0 626000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_393
timestamp 1765232829
transform 1 0 628000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_394
timestamp 1765232829
transform 1 0 699400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_396
timestamp 1765232829
transform 1 0 647800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_397
timestamp 1765232829
transform 1 0 649800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_398
timestamp 1765232829
transform 1 0 651800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_399
timestamp 1765232829
transform 1 0 653800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_402
timestamp 1765232829
transform 1 0 673600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_403
timestamp 1765232829
transform 1 0 675600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_404
timestamp 1765232829
transform 1 0 677600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_405
timestamp 1765232829
transform 1 0 679600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_406
timestamp 1765232829
transform 1 0 600200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_407
timestamp 1765232829
transform 1 0 594200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_408
timestamp 1765232829
transform 1 0 596200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_409
timestamp 1765232829
transform 1 0 598200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_410
timestamp 1765232829
transform 0 1 5200 -1 0 254500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_411
timestamp 1765232829
transform 1 0 391800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_412
timestamp 1765232829
transform 0 -1 781200 1 0 252500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_413
timestamp 1765232829
transform 1 0 391800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_0
timestamp 1765487709
transform 0 -1 781200 1 0 218300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_13
timestamp 1765487709
transform 1 0 671600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_22
timestamp 1765487709
transform 1 0 620000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_25
timestamp 1765487709
transform 1 0 645800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_36
timestamp 1765487709
transform 1 0 697400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_47
timestamp 1765487709
transform 1 0 465200 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_54
timestamp 1765487709
transform 1 0 491000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_58
timestamp 1765487709
transform 1 0 413600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_59
timestamp 1765487709
transform 1 0 542600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_65
timestamp 1765487709
transform 1 0 439400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_71
timestamp 1765487709
transform 1 0 516800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_78
timestamp 1765487709
transform 0 -1 781200 1 0 161900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_94
timestamp 1765487709
transform 0 -1 781200 1 0 246500
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_102
timestamp 1765487709
transform 0 -1 781200 1 0 190100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_103
timestamp 1765487709
transform 1 0 310400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_106
timestamp 1765487709
transform 1 0 258800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_113
timestamp 1765487709
transform 1 0 284600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_121
timestamp 1765487709
transform 1 0 336200 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_126
timestamp 1765487709
transform 1 0 362000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_138
timestamp 1765487709
transform 1 0 387800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_154
timestamp 1765487709
transform 1 0 104000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_163
timestamp 1765487709
transform 1 0 155600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_171
timestamp 1765487709
transform 1 0 181400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_177
timestamp 1765487709
transform 1 0 129800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_190
timestamp 1765487709
transform 0 1 5200 1 0 161900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_197
timestamp 1765487709
transform 0 1 5200 1 0 218300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_204
timestamp 1765487709
transform 0 1 5200 1 0 246500
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_205
timestamp 1765487709
transform 0 1 5200 1 0 190100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_247
timestamp 1765487709
transform 1 0 129800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_258
timestamp 1765487709
transform 1 0 181400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_264
timestamp 1765487709
transform 1 0 155600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_266
timestamp 1765487709
transform 1 0 104000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_271
timestamp 1765487709
transform 1 0 387800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_280
timestamp 1765487709
transform 1 0 284600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_287
timestamp 1765487709
transform 1 0 362000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_294
timestamp 1765487709
transform 1 0 310400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_300
timestamp 1765487709
transform 1 0 258800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_307
timestamp 1765487709
transform 1 0 336200 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_318
timestamp 1765487709
transform 0 -1 781200 1 0 274700
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_323
timestamp 1765487709
transform 0 -1 781200 1 0 359300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_331
timestamp 1765487709
transform 0 -1 781200 1 0 331100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_336
timestamp 1765487709
transform 1 0 413600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_341
timestamp 1765487709
transform 1 0 439400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_345
timestamp 1765487709
transform 1 0 465200 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_350
timestamp 1765487709
transform 1 0 491000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_355
timestamp 1765487709
transform 1 0 516800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_361
timestamp 1765487709
transform 1 0 542600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_389
timestamp 1765487709
transform 1 0 620000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_395
timestamp 1765487709
transform 1 0 645800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_400
timestamp 1765487709
transform 1 0 697400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_401
timestamp 1765487709
transform 1 0 671600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 90460
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_1
timestamp 1765232829
transform 0 -1 781200 1 0 90480
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_2
timestamp 1765232829
transform 0 -1 781200 1 0 90400
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_3
timestamp 1765232829
transform 0 -1 781200 1 0 90420
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_4
timestamp 1765232829
transform 0 -1 781200 1 0 90440
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_5
timestamp 1765232829
transform 0 1 5200 -1 0 90480
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_6
timestamp 1765232829
transform 0 1 5200 -1 0 90440
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_7
timestamp 1765232829
transform 0 1 5200 -1 0 90420
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_8
timestamp 1765232829
transform 0 1 5200 -1 0 90460
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_9
timestamp 1765232829
transform 0 1 5200 -1 0 90500
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_10
timestamp 1765232829
transform 0 1 5200 -1 0 430000
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_11
timestamp 1765232829
transform 0 1 5200 -1 0 429920
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_12
timestamp 1765232829
transform 0 1 5200 -1 0 429940
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_13
timestamp 1765232829
transform 0 1 5200 -1 0 429960
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_14
timestamp 1765232829
transform 0 1 5200 -1 0 429980
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_15
timestamp 1765232829
transform 0 -1 781200 1 0 429900
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_16
timestamp 1765232829
transform 0 -1 781200 1 0 429920
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_17
timestamp 1765232829
transform 0 -1 781200 1 0 429940
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_18
timestamp 1765232829
transform 0 -1 781200 1 0 429960
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_19
timestamp 1765232829
transform 0 -1 781200 1 0 429980
box -32 13097 52 69968
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform -1 0 129800 0 1 5200
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_1
timestamp 1765232829
transform 0 1 5200 -1 0 161900
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_2
timestamp 1765232829
transform 0 1 5200 -1 0 190100
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_3
timestamp 1765232829
transform 0 1 5200 -1 0 218300
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_4
timestamp 1765232829
transform 0 1 5200 -1 0 246500
box -32 0 15032 69970
use gf180mcu_ocd_io__in_s  gf180mcu_ocd_io__in_s_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform -1 0 104000 0 1 5200
box -32 0 15032 69970
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 118700
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_2
timestamp 1765232829
transform 1 0 218000 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_4
timestamp 1765232829
transform 0 1 5200 -1 0 415700
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_7
timestamp 1765232829
transform 1 0 579200 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765232829
transform 0 -1 781200 1 0 90500
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_3
timestamp 1765232829
transform 1 0 192200 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_4
timestamp 1765232829
transform 0 1 5200 -1 0 387500
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_6
timestamp 1765232829
transform 1 0 553400 0 -1 501000
box -32 0 15032 70000
use horz_connects  horz_connects_0
timestamp 1765054368
transform 1 0 141090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_1
timestamp 1765054368
transform 1 0 166890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_2
timestamp 1765054368
transform 1 0 244290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_3
timestamp 1765054368
transform 1 0 270090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_4
timestamp 1765054368
transform 1 0 295890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_5
timestamp 1765054368
transform 1 0 321690 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_6
timestamp 1765054368
transform 1 0 347490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_7
timestamp 1765054368
transform 1 0 373290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_8
timestamp 1765054368
transform 1 0 399090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_9
timestamp 1765054368
transform 1 0 424890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_10
timestamp 1765054368
transform 1 0 450690 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_11
timestamp 1765054368
transform 1 0 476490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_12
timestamp 1765054368
transform 1 0 502290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_13
timestamp 1765054368
transform 1 0 528090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_14
timestamp 1765054368
transform 1 0 605490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_15
timestamp 1765054368
transform 1 0 631290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_16
timestamp 1765054368
transform 1 0 657090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_17
timestamp 1765054368
transform 1 0 682890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_18
timestamp 1765054368
transform 1 0 682890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_19
timestamp 1765054368
transform 1 0 657090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_20
timestamp 1765054368
transform 1 0 631290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_21
timestamp 1765054368
transform 1 0 605490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_22
timestamp 1765054368
transform 1 0 528090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_23
timestamp 1765054368
transform 1 0 502290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_24
timestamp 1765054368
transform 1 0 476490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_25
timestamp 1765054368
transform 1 0 450690 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_26
timestamp 1765054368
transform 1 0 424890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_27
timestamp 1765054368
transform 1 0 399090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_28
timestamp 1765054368
transform 1 0 373290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_29
timestamp 1765054368
transform 1 0 347490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_30
timestamp 1765054368
transform 1 0 321690 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_31
timestamp 1765054368
transform 1 0 295890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_32
timestamp 1765054368
transform 1 0 270090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_33
timestamp 1765054368
transform 1 0 244290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_34
timestamp 1765054368
transform 1 0 166890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_35
timestamp 1765054368
transform 1 0 141090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_36
timestamp 1765054368
transform 1 0 115290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_37
timestamp 1765054368
transform 1 0 89490 0 -1 431000
box 0 -48 15527 232
use horz_connects_resetb  horz_connects_resetb_0
timestamp 1764982896
transform 1 0 115290 0 1 75170
box 12323 0 15527 232
use horz_connects_resetb  horz_connects_resetb_1
timestamp 1764982896
transform 1 0 89490 0 1 75170
box 12323 0 15527 232
use horz_power_connect  horz_power_connect_0
timestamp 1764102312
transform 1 0 192472 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_1
timestamp 1764102312
transform 1 0 218272 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_2
timestamp 1764102312
transform 1 0 553672 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_3
timestamp 1764102312
transform 1 0 579472 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_4
timestamp 1764102312
transform -1 0 593928 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_5
timestamp 1764102312
transform -1 0 568128 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_6
timestamp 1764102312
transform -1 0 232728 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_7
timestamp 1764102312
transform -1 0 206928 0 -1 431000
box 0 0 14456 200
use vert_connects  vert_connects_0
timestamp 1765055688
transform -1 0 711200 0 -1 162842
box 0 -67 303 15285
use vert_connects  vert_connects_1
timestamp 1765055688
transform -1 0 711200 0 -1 191042
box 0 -67 303 15285
use vert_connects  vert_connects_2
timestamp 1765055688
transform -1 0 711200 0 -1 219242
box 0 -67 303 15285
use vert_connects  vert_connects_3
timestamp 1765055688
transform -1 0 711200 0 -1 247442
box 0 -67 303 15285
use vert_connects  vert_connects_4
timestamp 1765055688
transform -1 0 711200 0 -1 275642
box 0 -67 303 15285
use vert_connects  vert_connects_5
timestamp 1765055688
transform -1 0 711200 0 -1 303842
box 0 -67 303 15285
use vert_connects  vert_connects_6
timestamp 1765055688
transform -1 0 711200 0 -1 332042
box 0 -67 303 15285
use vert_connects  vert_connects_7
timestamp 1765055688
transform -1 0 711200 0 -1 360242
box 0 -67 303 15285
use vert_connects_in_c  vert_connects_in_c_0
timestamp 1765055688
transform 1 0 75200 0 -1 191042
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_1
timestamp 1765055688
transform 1 0 75200 0 -1 162842
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_2
timestamp 1765055688
transform 1 0 75200 0 -1 219242
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_3
timestamp 1765055688
transform 1 0 75200 0 -1 247442
box -30 -62 303 15190
use vert_power_connect  vert_power_connect_0
timestamp 1764982451
transform 1 0 710930 0 1 90772
box 0 0 270 14456
use vert_power_connect  vert_power_connect_1
timestamp 1764982451
transform 1 0 710930 0 1 118972
box 0 0 270 14456
use vert_power_connect  vert_power_connect_2
timestamp 1764982451
transform 1 0 710930 0 1 372772
box 0 0 270 14456
use vert_power_connect  vert_power_connect_3
timestamp 1764982451
transform 1 0 710930 0 1 400972
box 0 0 270 14456
use vert_power_connect  vert_power_connect_4
timestamp 1764982451
transform -1 0 75470 0 -1 415428
box 0 0 270 14456
use vert_power_connect  vert_power_connect_5
timestamp 1764982451
transform -1 0 75470 0 -1 387228
box 0 0 270 14456
use vert_power_connect  vert_power_connect_6
timestamp 1764982451
transform -1 0 75470 0 -1 133428
box 0 0 270 14456
use vert_power_connect  vert_power_connect_7
timestamp 1764982451
transform -1 0 75470 0 -1 105228
box 0 0 270 14456
<< labels >>
rlabel metal5 s 584232 9168 589232 14168 4 DVDD
port 1 nsew
rlabel metal5 s 223032 9168 228032 14168 4 VDD
port 3 nsew
rlabel metal5 s 558432 9168 563432 14168 4 DVSS
port 2 nsew
rlabel metal5 s 197232 9168 202232 14168 4 VSS
port 4 nsew
rlabel metal5 s 584232 491968 589232 496968 4 VDD
port 3 nsew
rlabel metal5 s 223032 491968 228032 496968 4 DVDD
port 1 nsew
rlabel metal5 s 558432 491968 563432 496968 4 VSS
port 4 nsew
rlabel metal5 s 197232 491968 202232 496968 4 DVSS
port 2 nsew
rlabel metal5 s 9200 405732 14200 410732 4 VDD
port 3 nsew
rlabel metal5 s 9200 123732 14200 128732 4 DVDD
port 1 nsew
rlabel metal5 s 9200 377532 14200 382532 4 VSS
port 4 nsew
rlabel metal5 s 9200 95532 14200 100532 4 DVSS
port 2 nsew
rlabel metal5 s 772168 405732 777168 410732 4 DVDD
port 1 nsew
rlabel metal5 s 772168 123732 777168 128732 4 VDD
port 3 nsew
rlabel metal5 s 772168 377532 777168 382532 4 DVSS
port 2 nsew
rlabel metal5 s 772168 95532 777168 100532 4 VSS
port 4 nsew
rlabel metal5 9200 349332 14200 354332 0 analog_PAD[0]
port 55 nsew
rlabel metal5 9200 321132 14200 326132 0 analog_PAD[1]
port 54 nsew
rlabel metal5 9200 292932 14200 297932 0 analog_PAD[2]
port 53 nsew
rlabel metal5 9200 264732 14200 269732 0 analog_PAD[3]
port 52 nsew
rlabel metal5 9200 236532 14200 241532 0 input_PAD[0]
port 60 nsew
rlabel metal5 9200 208332 14200 213332 0 input_PAD[1]
port 59 nsew
rlabel metal5 9200 180132 14200 185132 0 input_PAD[2]
port 58 nsew
rlabel metal5 9200 151932 14200 156932 0 input_PAD[3]
port 57 nsew
rlabel metal5 94032 9168 99032 14168 0 clk_PAD
port 61 nsew
rlabel metal5 119832 9168 124832 14168 0 rst_n_PAD
port 62 nsew
rlabel metal5 145632 9168 150632 14168 0 bidir_PAD[0]
port 50 nsew
rlabel metal5 171432 9168 176432 14168 0 bidir_PAD[1]
port 49 nsew
rlabel metal5 248832 9168 253832 14168 0 bidir_PAD[2]
port 48 nsew
rlabel metal5 274632 9168 279632 14168 0 bidir_PAD[3]
port 47 nsew
rlabel metal5 300432 9168 305432 14168 0 bidir_PAD[4]
port 46 nsew
rlabel metal5 326232 9168 331232 14168 0 bidir_PAD[5]
port 45 nsew
rlabel metal5 352032 9168 357032 14168 0 bidir_PAD[6]
port 44 nsew
rlabel metal5 377832 9168 382832 14168 0 bidir_PAD[7]
port 43 nsew
rlabel metal5 403632 9168 408632 14168 0 bidir_PAD[8]
port 42 nsew
rlabel metal5 429432 9168 434432 14168 0 bidir_PAD[9]
port 41 nsew
rlabel metal5 455232 9168 460232 14168 0 bidir_PAD[10]
port 40 nsew
rlabel metal5 481032 9168 486032 14168 0 bidir_PAD[11]
port 39 nsew
rlabel metal5 506832 9168 511832 14168 0 bidir_PAD[12]
port 38 nsew
rlabel metal5 532632 9168 537632 14168 0 bidir_PAD[13]
port 37 nsew
rlabel metal5 610032 9168 615032 14168 0 bidir_PAD[14]
port 36 nsew
rlabel metal5 635832 9168 640832 14168 0 bidir_PAD[15]
port 35 nsew
rlabel metal5 661632 9168 666632 14168 0 bidir_PAD[16]
port 34 nsew
rlabel metal5 687432 9168 692432 14168 0 bidir_PAD[17]
port 33 nsew
rlabel metal5 772168 151932 777168 156932 0 bidir_PAD[18]
port 32 nsew
rlabel metal5 772168 180132 777168 185132 0 bidir_PAD[19]
port 31 nsew
rlabel metal5 772168 208332 777168 213332 0 bidir_PAD[20]
port 30 nsew
rlabel metal5 772168 236532 777168 241532 0 bidir_PAD[21]
port 29 nsew
rlabel metal5 772168 264732 777168 269732 0 bidir_PAD[22]
port 28 nsew
rlabel metal5 772168 292932 777168 297932 0 bidir_PAD[23]
port 27 nsew
rlabel metal5 772168 321132 777168 326132 0 bidir_PAD[24]
port 26 nsew
rlabel metal5 772168 349332 777168 354332 0 bidir_PAD[25]
port 25 nsew
rlabel metal5 687432 491968 692432 496968 0 bidir_PAD[26]
port 24 nsew
rlabel metal5 661632 491968 666632 496968 0 bidir_PAD[27]
port 23 nsew
rlabel metal5 635832 491968 640832 496968 0 bidir_PAD[28]
port 22 nsew
rlabel metal5 610032 491968 615032 496968 0 bidir_PAD[29]
port 21 nsew
rlabel metal5 532632 491968 537632 496968 0 bidir_PAD[30]
port 20 nsew
rlabel metal5 506832 491968 511832 496968 0 bidir_PAD[31]
port 19 nsew
rlabel metal5 481032 491968 486032 496968 0 bidir_PAD[32]
port 18 nsew
rlabel metal5 455232 491968 460232 496968 0 bidir_PAD[33]
port 17 nsew
rlabel metal5 429432 491968 434432 496968 0 bidir_PAD[34]
port 16 nsew
rlabel metal5 403632 491968 408632 496968 0 bidir_PAD[35]
port 15 nsew
rlabel metal5 377832 491968 382832 496968 0 bidir_PAD[36]
port 14 nsew
rlabel metal5 352032 491968 357032 496968 0 bidir_PAD[37]
port 13 nsew
rlabel metal5 326232 491968 331232 496968 0 bidir_PAD[38]
port 12 nsew
rlabel metal5 300432 491968 305432 496968 0 bidir_PAD[39]
port 11 nsew
rlabel metal5 274632 491968 279632 496968 0 bidir_PAD[40]
port 10 nsew
rlabel metal5 248832 491968 253832 496968 0 bidir_PAD[41]
port 9 nsew
rlabel metal5 171432 491968 176432 496968 0 bidir_PAD[42]
port 8 nsew
rlabel metal5 145632 491968 150632 496968 0 bidir_PAD[43]
port 7 nsew
rlabel metal5 119832 491968 124832 496968 0 bidir_PAD[44]
port 6 nsew
rlabel metal5 94032 491968 99032 496968 0 bidir_PAD[45]
port 5 nsew
flabel metal2 130546 75102 130622 75402 0 FreeSans 480 90 0 0 loopback_zero[51]
port 621 nsew
flabel metal2 130358 75102 130434 75402 0 FreeSans 480 90 0 0 loopback_one[51]
port 569 nsew
flabel metal2 128530 75102 128606 75402 0 FreeSans 480 90 0 0 rst_n_PU
port 691 nsew
flabel metal2 127658 75102 127734 75402 0 FreeSans 480 90 0 0 rst_n_PD
port 692 nsew
flabel metal2 104746 75102 104822 75402 0 FreeSans 480 90 0 0 loopback_zero[50]
port 622 nsew
flabel metal2 104558 75102 104634 75402 0 FreeSans 480 90 0 0 loopback_one[50]
port 570 nsew
flabel metal2 102730 75102 102806 75402 0 FreeSans 480 90 0 0 clk_PU
port 688 nsew
flabel metal2 101858 75102 101934 75402 0 FreeSans 480 90 0 0 clk_PD
port 689 nsew
flabel metal2 89752 75102 89826 75402 0 FreeSans 480 90 0 0 clk_Y
port 690 nsew
flabel metal2 115552 75102 115626 75402 0 FreeSans 480 90 0 0 rst_n_Y
port 693 nsew
flabel metal2 141272 75132 141348 75432 0 FreeSans 480 90 0 0 bidir_CS[0]
port 108 nsew
flabel metal2 141793 75132 141869 75432 0 FreeSans 480 90 0 0 bidir_PU[0]
port 154 nsew
flabel metal2 142022 75132 142098 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[0]
port 200 nsew
flabel metal2 142164 75132 142240 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[0]
port 246 nsew
flabel metal2 142666 75132 142742 75432 0 FreeSans 480 90 0 0 bidir_PD[0]
port 338 nsew
flabel metal2 142877 75132 142953 75432 0 FreeSans 480 90 0 0 bidir_IE[0]
port 384 nsew
flabel metal2 142306 75132 142382 75432 0 FreeSans 480 90 0 0 bidir_ANA[0]
port 292 nsew
flabel metal2 154334 75132 154410 75432 0 FreeSans 480 90 0 0 bidir_SL[0]
port 430 nsew
flabel metal2 154480 75132 154556 75432 0 FreeSans 480 90 0 0 bidir_A[0]
port 476 nsew
flabel metal2 154626 75132 154702 75432 0 FreeSans 480 90 0 0 bidir_OE[0]
port 522 nsew
flabel metal2 154772 75132 154848 75432 0 FreeSans 480 90 0 0 bidir_Y[0]
port 568 nsew
flabel metal2 156158 75132 156234 75432 0 FreeSans 480 90 0 0 loopback_one[0]
port 620 nsew
flabel metal2 156346 75132 156422 75432 0 FreeSans 480 90 0 0 loopback_zero[0]
port 672 nsew
flabel metal2 167072 75132 167148 75432 0 FreeSans 480 90 0 0 bidir_CS[1]
port 107 nsew
flabel metal2 167593 75132 167669 75432 0 FreeSans 480 90 0 0 bidir_PU[1]
port 153 nsew
flabel metal2 167822 75132 167898 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[1]
port 199 nsew
flabel metal2 167964 75132 168040 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[1]
port 245 nsew
flabel metal2 168106 75132 168182 75432 0 FreeSans 480 90 0 0 bidir_ANA[1]
port 291 nsew
flabel metal2 168466 75132 168542 75432 0 FreeSans 480 90 0 0 bidir_PD[1]
port 337 nsew
flabel metal2 168677 75132 168753 75432 0 FreeSans 480 90 0 0 bidir_IE[1]
port 383 nsew
flabel metal2 180134 75132 180210 75432 0 FreeSans 480 90 0 0 bidir_SL[1]
port 429 nsew
flabel metal2 180280 75132 180356 75432 0 FreeSans 480 90 0 0 bidir_A[1]
port 475 nsew
flabel metal2 180426 75132 180502 75432 0 FreeSans 480 90 0 0 bidir_OE[1]
port 521 nsew
flabel metal2 180572 75132 180648 75432 0 FreeSans 480 90 0 0 bidir_Y[1]
port 567 nsew
flabel metal2 181958 75132 182034 75432 0 FreeSans 480 90 0 0 loopback_one[1]
port 619 nsew
flabel metal2 182146 75132 182222 75432 0 FreeSans 480 90 0 0 loopback_zero[1]
port 671 nsew
flabel metal2 259546 75132 259622 75432 0 FreeSans 480 90 0 0 loopback_zero[2]
port 670 nsew
flabel metal2 259358 75132 259434 75432 0 FreeSans 480 90 0 0 loopback_one[2]
port 618 nsew
flabel metal2 257972 75132 258048 75432 0 FreeSans 480 90 0 0 bidir_Y[2]
port 566 nsew
flabel metal2 257826 75132 257902 75432 0 FreeSans 480 90 0 0 bidir_OE[2]
port 520 nsew
flabel metal2 257680 75132 257756 75432 0 FreeSans 480 90 0 0 bidir_A[2]
port 474 nsew
flabel metal2 257534 75132 257610 75432 0 FreeSans 480 90 0 0 bidir_SL[2]
port 428 nsew
flabel metal2 246077 75132 246153 75432 0 FreeSans 480 90 0 0 bidir_IE[2]
port 382 nsew
flabel metal2 245866 75132 245942 75432 0 FreeSans 480 90 0 0 bidir_PD[2]
port 336 nsew
flabel metal2 245506 75132 245582 75432 0 FreeSans 480 90 0 0 bidir_ANA[2]
port 290 nsew
flabel metal2 245364 75132 245440 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[2]
port 244 nsew
flabel metal2 245222 75132 245298 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[2]
port 198 nsew
flabel metal2 244993 75132 245069 75432 0 FreeSans 480 90 0 0 bidir_PU[2]
port 152 nsew
flabel metal2 244472 75132 244548 75432 0 FreeSans 480 90 0 0 bidir_CS[2]
port 106 nsew
flabel metal2 285346 75132 285422 75432 0 FreeSans 480 90 0 0 loopback_zero[3]
port 669 nsew
flabel metal2 285158 75132 285234 75432 0 FreeSans 480 90 0 0 loopback_one[3]
port 617 nsew
flabel metal2 283772 75132 283848 75432 0 FreeSans 480 90 0 0 bidir_Y[3]
port 565 nsew
flabel metal2 283626 75132 283702 75432 0 FreeSans 480 90 0 0 bidir_OE[3]
port 519 nsew
flabel metal2 283480 75132 283556 75432 0 FreeSans 480 90 0 0 bidir_A[3]
port 473 nsew
flabel metal2 283334 75132 283410 75432 0 FreeSans 480 90 0 0 bidir_SL[3]
port 427 nsew
flabel metal2 271877 75132 271953 75432 0 FreeSans 480 90 0 0 bidir_IE[3]
port 381 nsew
flabel metal2 271666 75132 271742 75432 0 FreeSans 480 90 0 0 bidir_PD[3]
port 335 nsew
flabel metal2 271306 75132 271382 75432 0 FreeSans 480 90 0 0 bidir_ANA[3]
port 289 nsew
flabel metal2 271164 75132 271240 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[3]
port 243 nsew
flabel metal2 271022 75132 271098 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[3]
port 197 nsew
flabel metal2 270793 75132 270869 75432 0 FreeSans 480 90 0 0 bidir_PU[3]
port 151 nsew
flabel metal2 270272 75132 270348 75432 0 FreeSans 480 90 0 0 bidir_CS[3]
port 105 nsew
flabel metal2 311146 75132 311222 75432 0 FreeSans 480 90 0 0 loopback_zero[4]
port 668 nsew
flabel metal2 310958 75132 311034 75432 0 FreeSans 480 90 0 0 loopback_one[4]
port 616 nsew
flabel metal2 309572 75132 309648 75432 0 FreeSans 480 90 0 0 bidir_Y[4]
port 564 nsew
flabel metal2 309426 75132 309502 75432 0 FreeSans 480 90 0 0 bidir_OE[4]
port 518 nsew
flabel metal2 309280 75132 309356 75432 0 FreeSans 480 90 0 0 bidir_A[4]
port 472 nsew
flabel metal2 309134 75132 309210 75432 0 FreeSans 480 90 0 0 bidir_SL[4]
port 426 nsew
flabel metal2 297677 75132 297753 75432 0 FreeSans 480 90 0 0 bidir_IE[4]
port 380 nsew
flabel metal2 297466 75132 297542 75432 0 FreeSans 480 90 0 0 bidir_PD[4]
port 334 nsew
flabel metal2 297106 75132 297182 75432 0 FreeSans 480 90 0 0 bidir_ANA[4]
port 288 nsew
flabel metal2 296964 75132 297040 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[4]
port 242 nsew
flabel metal2 296822 75132 296898 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[4]
port 196 nsew
flabel metal2 296593 75132 296669 75432 0 FreeSans 480 90 0 0 bidir_PU[4]
port 150 nsew
flabel metal2 296072 75132 296148 75432 0 FreeSans 480 90 0 0 bidir_CS[4]
port 104 nsew
flabel metal2 336946 75132 337022 75432 0 FreeSans 480 90 0 0 loopback_zero[5]
port 667 nsew
flabel metal2 336758 75132 336834 75432 0 FreeSans 480 90 0 0 loopback_one[5]
port 615 nsew
flabel metal2 335372 75132 335448 75432 0 FreeSans 480 90 0 0 bidir_Y[5]
port 563 nsew
flabel metal2 335226 75132 335302 75432 0 FreeSans 480 90 0 0 bidir_OE[5]
port 517 nsew
flabel metal2 335080 75132 335156 75432 0 FreeSans 480 90 0 0 bidir_A[5]
port 471 nsew
flabel metal2 334934 75132 335010 75432 0 FreeSans 480 90 0 0 bidir_SL[5]
port 425 nsew
flabel metal2 323477 75132 323553 75432 0 FreeSans 480 90 0 0 bidir_IE[5]
port 379 nsew
flabel metal2 323266 75132 323342 75432 0 FreeSans 480 90 0 0 bidir_PD[5]
port 333 nsew
flabel metal2 322906 75132 322982 75432 0 FreeSans 480 90 0 0 bidir_ANA[5]
port 287 nsew
flabel metal2 322764 75132 322840 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[5]
port 241 nsew
flabel metal2 322622 75132 322698 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[5]
port 195 nsew
flabel metal2 322393 75132 322469 75432 0 FreeSans 480 90 0 0 bidir_PU[5]
port 149 nsew
flabel metal2 321872 75132 321948 75432 0 FreeSans 480 90 0 0 bidir_CS[5]
port 103 nsew
flabel metal2 362746 75132 362822 75432 0 FreeSans 480 90 0 0 loopback_zero[6]
port 666 nsew
flabel metal2 362558 75132 362634 75432 0 FreeSans 480 90 0 0 loopback_one[6]
port 614 nsew
flabel metal2 361172 75132 361248 75432 0 FreeSans 480 90 0 0 bidir_Y[6]
port 562 nsew
flabel metal2 361026 75132 361102 75432 0 FreeSans 480 90 0 0 bidir_OE[6]
port 516 nsew
flabel metal2 360880 75132 360956 75432 0 FreeSans 480 90 0 0 bidir_A[6]
port 470 nsew
flabel metal2 360734 75132 360810 75432 0 FreeSans 480 90 0 0 bidir_SL[6]
port 424 nsew
flabel metal2 349277 75132 349353 75432 0 FreeSans 480 90 0 0 bidir_IE[6]
port 378 nsew
flabel metal2 349066 75132 349142 75432 0 FreeSans 480 90 0 0 bidir_PD[6]
port 332 nsew
flabel metal2 348706 75132 348782 75432 0 FreeSans 480 90 0 0 bidir_ANA[6]
port 286 nsew
flabel metal2 348564 75132 348640 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[6]
port 240 nsew
flabel metal2 348422 75132 348498 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[6]
port 194 nsew
flabel metal2 348193 75132 348269 75432 0 FreeSans 480 90 0 0 bidir_PU[6]
port 148 nsew
flabel metal2 347672 75132 347748 75432 0 FreeSans 480 90 0 0 bidir_CS[6]
port 102 nsew
flabel metal2 388546 75132 388622 75432 0 FreeSans 480 90 0 0 loopback_zero[7]
port 665 nsew
flabel metal2 388358 75132 388434 75432 0 FreeSans 480 90 0 0 loopback_one[7]
port 613 nsew
flabel metal2 386972 75132 387048 75432 0 FreeSans 480 90 0 0 bidir_Y[7]
port 561 nsew
flabel metal2 386826 75132 386902 75432 0 FreeSans 480 90 0 0 bidir_OE[7]
port 515 nsew
flabel metal2 386680 75132 386756 75432 0 FreeSans 480 90 0 0 bidir_A[7]
port 469 nsew
flabel metal2 386534 75132 386610 75432 0 FreeSans 480 90 0 0 bidir_SL[7]
port 423 nsew
flabel metal2 375077 75132 375153 75432 0 FreeSans 480 90 0 0 bidir_IE[7]
port 377 nsew
flabel metal2 374866 75132 374942 75432 0 FreeSans 480 90 0 0 bidir_PD[7]
port 331 nsew
flabel metal2 374506 75132 374582 75432 0 FreeSans 480 90 0 0 bidir_ANA[7]
port 285 nsew
flabel metal2 374364 75132 374440 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[7]
port 239 nsew
flabel metal2 374222 75132 374298 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[7]
port 193 nsew
flabel metal2 373993 75132 374069 75432 0 FreeSans 480 90 0 0 bidir_PU[7]
port 147 nsew
flabel metal2 373472 75132 373548 75432 0 FreeSans 480 90 0 0 bidir_CS[7]
port 101 nsew
flabel metal2 414346 75132 414422 75432 0 FreeSans 480 90 0 0 loopback_zero[8]
port 664 nsew
flabel metal2 414158 75132 414234 75432 0 FreeSans 480 90 0 0 loopback_one[8]
port 612 nsew
flabel metal2 412772 75132 412848 75432 0 FreeSans 480 90 0 0 bidir_Y[8]
port 560 nsew
flabel metal2 412626 75132 412702 75432 0 FreeSans 480 90 0 0 bidir_OE[8]
port 514 nsew
flabel metal2 412480 75132 412556 75432 0 FreeSans 480 90 0 0 bidir_A[8]
port 468 nsew
flabel metal2 412334 75132 412410 75432 0 FreeSans 480 90 0 0 bidir_SL[8]
port 422 nsew
flabel metal2 400877 75132 400953 75432 0 FreeSans 480 90 0 0 bidir_IE[8]
port 376 nsew
flabel metal2 400666 75132 400742 75432 0 FreeSans 480 90 0 0 bidir_PD[8]
port 330 nsew
flabel metal2 400306 75132 400382 75432 0 FreeSans 480 90 0 0 bidir_ANA[8]
port 284 nsew
flabel metal2 400164 75132 400240 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[8]
port 238 nsew
flabel metal2 400022 75132 400098 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[8]
port 192 nsew
flabel metal2 399793 75132 399869 75432 0 FreeSans 480 90 0 0 bidir_PU[8]
port 146 nsew
flabel metal2 399272 75132 399348 75432 0 FreeSans 480 90 0 0 bidir_CS[8]
port 100 nsew
flabel metal2 440146 75132 440222 75432 0 FreeSans 480 90 0 0 loopback_zero[9]
port 663 nsew
flabel metal2 439958 75132 440034 75432 0 FreeSans 480 90 0 0 loopback_one[9]
port 611 nsew
flabel metal2 438572 75132 438648 75432 0 FreeSans 480 90 0 0 bidir_Y[9]
port 559 nsew
flabel metal2 438426 75132 438502 75432 0 FreeSans 480 90 0 0 bidir_OE[9]
port 513 nsew
flabel metal2 438280 75132 438356 75432 0 FreeSans 480 90 0 0 bidir_A[9]
port 467 nsew
flabel metal2 438134 75132 438210 75432 0 FreeSans 480 90 0 0 bidir_SL[9]
port 421 nsew
flabel metal2 426677 75132 426753 75432 0 FreeSans 480 90 0 0 bidir_IE[9]
port 375 nsew
flabel metal2 426466 75132 426542 75432 0 FreeSans 480 90 0 0 bidir_PD[9]
port 329 nsew
flabel metal2 426106 75132 426182 75432 0 FreeSans 480 90 0 0 bidir_ANA[9]
port 283 nsew
flabel metal2 425964 75132 426040 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[9]
port 237 nsew
flabel metal2 425822 75132 425898 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[9]
port 191 nsew
flabel metal2 425593 75132 425669 75432 0 FreeSans 480 90 0 0 bidir_PU[9]
port 145 nsew
flabel metal2 425072 75132 425148 75432 0 FreeSans 480 90 0 0 bidir_CS[9]
port 99 nsew
flabel metal2 465946 75132 466022 75432 0 FreeSans 480 90 0 0 loopback_zero[10]
port 662 nsew
flabel metal2 465758 75132 465834 75432 0 FreeSans 480 90 0 0 loopback_one[10]
port 610 nsew
flabel metal2 464372 75132 464448 75432 0 FreeSans 480 90 0 0 bidir_Y[10]
port 558 nsew
flabel metal2 464226 75132 464302 75432 0 FreeSans 480 90 0 0 bidir_OE[10]
port 512 nsew
flabel metal2 464080 75132 464156 75432 0 FreeSans 480 90 0 0 bidir_A[10]
port 466 nsew
flabel metal2 463934 75132 464010 75432 0 FreeSans 480 90 0 0 bidir_SL[10]
port 420 nsew
flabel metal2 452477 75132 452553 75432 0 FreeSans 480 90 0 0 bidir_IE[10]
port 374 nsew
flabel metal2 452266 75132 452342 75432 0 FreeSans 480 90 0 0 bidir_PD[10]
port 328 nsew
flabel metal2 451906 75132 451982 75432 0 FreeSans 480 90 0 0 bidir_ANA[10]
port 282 nsew
flabel metal2 451764 75132 451840 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[10]
port 236 nsew
flabel metal2 451622 75132 451698 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[10]
port 190 nsew
flabel metal2 451393 75132 451469 75432 0 FreeSans 480 90 0 0 bidir_PU[10]
port 144 nsew
flabel metal2 450872 75132 450948 75432 0 FreeSans 480 90 0 0 bidir_CS[10]
port 98 nsew
flabel metal2 491746 75132 491822 75432 0 FreeSans 480 90 0 0 loopback_zero[11]
port 661 nsew
flabel metal2 491558 75132 491634 75432 0 FreeSans 480 90 0 0 loopback_one[11]
port 609 nsew
flabel metal2 490172 75132 490248 75432 0 FreeSans 480 90 0 0 bidir_Y[11]
port 557 nsew
flabel metal2 490026 75132 490102 75432 0 FreeSans 480 90 0 0 bidir_OE[11]
port 511 nsew
flabel metal2 489880 75132 489956 75432 0 FreeSans 480 90 0 0 bidir_A[11]
port 465 nsew
flabel metal2 489734 75132 489810 75432 0 FreeSans 480 90 0 0 bidir_SL[11]
port 419 nsew
flabel metal2 478277 75132 478353 75432 0 FreeSans 480 90 0 0 bidir_IE[11]
port 373 nsew
flabel metal2 478066 75132 478142 75432 0 FreeSans 480 90 0 0 bidir_PD[11]
port 327 nsew
flabel metal2 477706 75132 477782 75432 0 FreeSans 480 90 0 0 bidir_ANA[11]
port 281 nsew
flabel metal2 477564 75132 477640 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[11]
port 235 nsew
flabel metal2 477422 75132 477498 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[11]
port 189 nsew
flabel metal2 477193 75132 477269 75432 0 FreeSans 480 90 0 0 bidir_PU[11]
port 143 nsew
flabel metal2 476672 75132 476748 75432 0 FreeSans 480 90 0 0 bidir_CS[11]
port 97 nsew
flabel metal2 517546 75132 517622 75432 0 FreeSans 480 90 0 0 loopback_zero[12]
port 660 nsew
flabel metal2 517358 75132 517434 75432 0 FreeSans 480 90 0 0 loopback_one[12]
port 608 nsew
flabel metal2 515972 75132 516048 75432 0 FreeSans 480 90 0 0 bidir_Y[12]
port 556 nsew
flabel metal2 515826 75132 515902 75432 0 FreeSans 480 90 0 0 bidir_OE[12]
port 510 nsew
flabel metal2 515680 75132 515756 75432 0 FreeSans 480 90 0 0 bidir_A[12]
port 464 nsew
flabel metal2 515534 75132 515610 75432 0 FreeSans 480 90 0 0 bidir_SL[12]
port 418 nsew
flabel metal2 504077 75132 504153 75432 0 FreeSans 480 90 0 0 bidir_IE[12]
port 372 nsew
flabel metal2 503866 75132 503942 75432 0 FreeSans 480 90 0 0 bidir_PD[12]
port 326 nsew
flabel metal2 503506 75132 503582 75432 0 FreeSans 480 90 0 0 bidir_ANA[12]
port 280 nsew
flabel metal2 503364 75132 503440 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[12]
port 234 nsew
flabel metal2 503222 75132 503298 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[12]
port 188 nsew
flabel metal2 502993 75132 503069 75432 0 FreeSans 480 90 0 0 bidir_PU[12]
port 142 nsew
flabel metal2 502472 75132 502548 75432 0 FreeSans 480 90 0 0 bidir_CS[12]
port 96 nsew
flabel metal2 543346 75132 543422 75432 0 FreeSans 480 90 0 0 loopback_zero[13]
port 659 nsew
flabel metal2 543158 75132 543234 75432 0 FreeSans 480 90 0 0 loopback_one[13]
port 607 nsew
flabel metal2 541772 75132 541848 75432 0 FreeSans 480 90 0 0 bidir_Y[13]
port 555 nsew
flabel metal2 541626 75132 541702 75432 0 FreeSans 480 90 0 0 bidir_OE[13]
port 509 nsew
flabel metal2 541480 75132 541556 75432 0 FreeSans 480 90 0 0 bidir_A[13]
port 463 nsew
flabel metal2 541334 75132 541410 75432 0 FreeSans 480 90 0 0 bidir_SL[13]
port 417 nsew
flabel metal2 529877 75132 529953 75432 0 FreeSans 480 90 0 0 bidir_IE[13]
port 371 nsew
flabel metal2 529666 75132 529742 75432 0 FreeSans 480 90 0 0 bidir_PD[13]
port 325 nsew
flabel metal2 529306 75132 529382 75432 0 FreeSans 480 90 0 0 bidir_ANA[13]
port 279 nsew
flabel metal2 529164 75132 529240 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[13]
port 233 nsew
flabel metal2 529022 75132 529098 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[13]
port 187 nsew
flabel metal2 528793 75132 528869 75432 0 FreeSans 480 90 0 0 bidir_PU[13]
port 141 nsew
flabel metal2 528272 75132 528348 75432 0 FreeSans 480 90 0 0 bidir_CS[13]
port 95 nsew
flabel metal2 620746 75132 620822 75432 0 FreeSans 480 90 0 0 loopback_zero[14]
port 658 nsew
flabel metal2 620558 75132 620634 75432 0 FreeSans 480 90 0 0 loopback_one[14]
port 606 nsew
flabel metal2 619172 75132 619248 75432 0 FreeSans 480 90 0 0 bidir_Y[14]
port 554 nsew
flabel metal2 619026 75132 619102 75432 0 FreeSans 480 90 0 0 bidir_OE[14]
port 508 nsew
flabel metal2 618880 75132 618956 75432 0 FreeSans 480 90 0 0 bidir_A[14]
port 462 nsew
flabel metal2 618734 75132 618810 75432 0 FreeSans 480 90 0 0 bidir_SL[14]
port 416 nsew
flabel metal2 607277 75132 607353 75432 0 FreeSans 480 90 0 0 bidir_IE[14]
port 370 nsew
flabel metal2 607066 75132 607142 75432 0 FreeSans 480 90 0 0 bidir_PD[14]
port 324 nsew
flabel metal2 606706 75132 606782 75432 0 FreeSans 480 90 0 0 bidir_ANA[14]
port 278 nsew
flabel metal2 606564 75132 606640 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[14]
port 232 nsew
flabel metal2 606422 75132 606498 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[14]
port 186 nsew
flabel metal2 606193 75132 606269 75432 0 FreeSans 480 90 0 0 bidir_PU[14]
port 140 nsew
flabel metal2 605672 75132 605748 75432 0 FreeSans 480 90 0 0 bidir_CS[14]
port 94 nsew
flabel metal2 646546 75132 646622 75432 0 FreeSans 480 90 0 0 loopback_zero[15]
port 657 nsew
flabel metal2 646358 75132 646434 75432 0 FreeSans 480 90 0 0 loopback_one[15]
port 605 nsew
flabel metal2 644972 75132 645048 75432 0 FreeSans 480 90 0 0 bidir_Y[15]
port 553 nsew
flabel metal2 644826 75132 644902 75432 0 FreeSans 480 90 0 0 bidir_OE[15]
port 507 nsew
flabel metal2 644680 75132 644756 75432 0 FreeSans 480 90 0 0 bidir_A[15]
port 461 nsew
flabel metal2 644534 75132 644610 75432 0 FreeSans 480 90 0 0 bidir_SL[15]
port 415 nsew
flabel metal2 633077 75132 633153 75432 0 FreeSans 480 90 0 0 bidir_IE[15]
port 369 nsew
flabel metal2 632866 75132 632942 75432 0 FreeSans 480 90 0 0 bidir_PD[15]
port 323 nsew
flabel metal2 632506 75132 632582 75432 0 FreeSans 480 90 0 0 bidir_ANA[15]
port 277 nsew
flabel metal2 632364 75132 632440 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[15]
port 231 nsew
flabel metal2 632222 75132 632298 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[15]
port 185 nsew
flabel metal2 631993 75132 632069 75432 0 FreeSans 480 90 0 0 bidir_PU[15]
port 139 nsew
flabel metal2 631472 75132 631548 75432 0 FreeSans 480 90 0 0 bidir_CS[15]
port 93 nsew
flabel metal2 672346 75132 672422 75432 0 FreeSans 480 90 0 0 loopback_zero[16]
port 656 nsew
flabel metal2 672158 75132 672234 75432 0 FreeSans 480 90 0 0 loopback_one[16]
port 604 nsew
flabel metal2 670772 75132 670848 75432 0 FreeSans 480 90 0 0 bidir_Y[16]
port 552 nsew
flabel metal2 670626 75132 670702 75432 0 FreeSans 480 90 0 0 bidir_OE[16]
port 506 nsew
flabel metal2 670480 75132 670556 75432 0 FreeSans 480 90 0 0 bidir_A[16]
port 460 nsew
flabel metal2 670334 75132 670410 75432 0 FreeSans 480 90 0 0 bidir_SL[16]
port 414 nsew
flabel metal2 658877 75132 658953 75432 0 FreeSans 480 90 0 0 bidir_IE[16]
port 368 nsew
flabel metal2 658666 75132 658742 75432 0 FreeSans 480 90 0 0 bidir_PD[16]
port 322 nsew
flabel metal2 658306 75132 658382 75432 0 FreeSans 480 90 0 0 bidir_ANA[16]
port 276 nsew
flabel metal2 658164 75132 658240 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[16]
port 230 nsew
flabel metal2 658022 75132 658098 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[16]
port 184 nsew
flabel metal2 657793 75132 657869 75432 0 FreeSans 480 90 0 0 bidir_PU[16]
port 138 nsew
flabel metal2 657272 75132 657348 75432 0 FreeSans 480 90 0 0 bidir_CS[16]
port 92 nsew
flabel metal2 698146 75132 698222 75432 0 FreeSans 480 90 0 0 loopback_zero[17]
port 655 nsew
flabel metal2 697958 75132 698034 75432 0 FreeSans 480 90 0 0 loopback_one[17]
port 603 nsew
flabel metal2 696572 75132 696648 75432 0 FreeSans 480 90 0 0 bidir_Y[17]
port 551 nsew
flabel metal2 696426 75132 696502 75432 0 FreeSans 480 90 0 0 bidir_OE[17]
port 505 nsew
flabel metal2 696280 75132 696356 75432 0 FreeSans 480 90 0 0 bidir_A[17]
port 459 nsew
flabel metal2 696134 75132 696210 75432 0 FreeSans 480 90 0 0 bidir_SL[17]
port 413 nsew
flabel metal2 684677 75132 684753 75432 0 FreeSans 480 90 0 0 bidir_IE[17]
port 367 nsew
flabel metal2 684466 75132 684542 75432 0 FreeSans 480 90 0 0 bidir_PD[17]
port 321 nsew
flabel metal2 684106 75132 684182 75432 0 FreeSans 480 90 0 0 bidir_ANA[17]
port 275 nsew
flabel metal2 683964 75132 684040 75432 0 FreeSans 480 90 0 0 bidir_PDRV1[17]
port 229 nsew
flabel metal2 683822 75132 683898 75432 0 FreeSans 480 90 0 0 bidir_PDRV0[17]
port 183 nsew
flabel metal2 683593 75132 683669 75432 0 FreeSans 480 90 0 0 bidir_PU[17]
port 137 nsew
flabel metal2 683072 75132 683148 75432 0 FreeSans 480 90 0 0 bidir_CS[17]
port 91 nsew
flabel metal3 710897 147572 711197 147648 0 FreeSans 480 0 0 0 bidir_CS[18]
port 90 nsew
flabel metal3 710897 148093 711197 148169 0 FreeSans 480 0 0 0 bidir_PU[18]
port 136 nsew
flabel metal3 710897 148322 711197 148398 0 FreeSans 480 0 0 0 bidir_PDRV0[18]
port 182 nsew
flabel metal3 710897 148464 711197 148540 0 FreeSans 480 0 0 0 bidir_PDRV1[18]
port 228 nsew
flabel metal3 710897 148606 711197 148682 0 FreeSans 480 0 0 0 bidir_ANA[18]
port 274 nsew
flabel metal3 710897 148966 711197 149042 0 FreeSans 480 0 0 0 bidir_PD[18]
port 320 nsew
flabel metal3 710897 149177 711197 149253 0 FreeSans 480 0 0 0 bidir_IE[18]
port 366 nsew
flabel metal3 710897 160634 711197 160710 0 FreeSans 480 0 0 0 bidir_SL[18]
port 412 nsew
flabel metal3 710897 160780 711197 160856 0 FreeSans 480 0 0 0 bidir_A[18]
port 458 nsew
flabel metal3 710897 160926 711197 161002 0 FreeSans 480 0 0 0 bidir_OE[18]
port 504 nsew
flabel metal3 710897 161072 711197 161148 0 FreeSans 480 0 0 0 bidir_Y[18]
port 550 nsew
flabel metal3 710897 162458 711197 162534 0 FreeSans 480 0 0 0 loopback_one[18]
port 602 nsew
flabel metal3 710897 162646 711197 162722 0 FreeSans 480 0 0 0 loopback_zero[18]
port 654 nsew
flabel metal3 710897 175772 711197 175848 0 FreeSans 480 0 0 0 bidir_CS[19]
port 89 nsew
flabel metal3 710897 176293 711197 176369 0 FreeSans 480 0 0 0 bidir_PU[19]
port 135 nsew
flabel metal3 710897 176522 711197 176598 0 FreeSans 480 0 0 0 bidir_PDRV0[19]
port 181 nsew
flabel metal3 710897 176664 711197 176740 0 FreeSans 480 0 0 0 bidir_PDRV1[19]
port 227 nsew
flabel metal3 710897 176806 711197 176882 0 FreeSans 480 0 0 0 bidir_ANA[19]
port 273 nsew
flabel metal3 710897 177166 711197 177242 0 FreeSans 480 0 0 0 bidir_PD[19]
port 319 nsew
flabel metal3 710897 177377 711197 177453 0 FreeSans 480 0 0 0 bidir_IE[19]
port 365 nsew
flabel metal3 710897 188834 711197 188910 0 FreeSans 480 0 0 0 bidir_SL[19]
port 411 nsew
flabel metal3 710897 188980 711197 189056 0 FreeSans 480 0 0 0 bidir_A[19]
port 457 nsew
flabel metal3 710897 189126 711197 189202 0 FreeSans 480 0 0 0 bidir_OE[19]
port 503 nsew
flabel metal3 710897 189272 711197 189348 0 FreeSans 480 0 0 0 bidir_Y[19]
port 549 nsew
flabel metal3 710897 190658 711197 190734 0 FreeSans 480 0 0 0 loopback_one[19]
port 601 nsew
flabel metal3 710897 190846 711197 190922 0 FreeSans 480 0 0 0 loopback_zero[19]
port 653 nsew
flabel metal3 710897 203972 711197 204048 0 FreeSans 480 0 0 0 bidir_CS[20]
port 88 nsew
flabel metal3 710897 204493 711197 204569 0 FreeSans 480 0 0 0 bidir_PU[20]
port 134 nsew
flabel metal3 710897 204722 711197 204798 0 FreeSans 480 0 0 0 bidir_PDRV0[20]
port 180 nsew
flabel metal3 710897 204864 711197 204940 0 FreeSans 480 0 0 0 bidir_PDRV1[20]
port 226 nsew
flabel metal3 710897 205006 711197 205082 0 FreeSans 480 0 0 0 bidir_ANA[20]
port 272 nsew
flabel metal3 710897 205366 711197 205442 0 FreeSans 480 0 0 0 bidir_PD[20]
port 318 nsew
flabel metal3 710897 205577 711197 205653 0 FreeSans 480 0 0 0 bidir_IE[20]
port 364 nsew
flabel metal3 710897 217034 711197 217110 0 FreeSans 480 0 0 0 bidir_SL[20]
port 410 nsew
flabel metal3 710897 217180 711197 217256 0 FreeSans 480 0 0 0 bidir_A[20]
port 456 nsew
flabel metal3 710897 217326 711197 217402 0 FreeSans 480 0 0 0 bidir_OE[20]
port 502 nsew
flabel metal3 710897 217472 711197 217548 0 FreeSans 480 0 0 0 bidir_Y[20]
port 548 nsew
flabel metal3 710897 218858 711197 218934 0 FreeSans 480 0 0 0 loopback_one[20]
port 600 nsew
flabel metal3 710897 219046 711197 219122 0 FreeSans 480 0 0 0 loopback_zero[20]
port 652 nsew
flabel metal3 710897 232172 711197 232248 0 FreeSans 480 0 0 0 bidir_CS[21]
port 87 nsew
flabel metal3 710897 232693 711197 232769 0 FreeSans 480 0 0 0 bidir_PU[21]
port 133 nsew
flabel metal3 710897 232922 711197 232998 0 FreeSans 480 0 0 0 bidir_PDRV0[21]
port 179 nsew
flabel metal3 710897 233064 711197 233140 0 FreeSans 480 0 0 0 bidir_PDRV1[21]
port 225 nsew
flabel metal3 710897 233206 711197 233282 0 FreeSans 480 0 0 0 bidir_ANA[21]
port 271 nsew
flabel metal3 710897 233566 711197 233642 0 FreeSans 480 0 0 0 bidir_PD[21]
port 317 nsew
flabel metal3 710897 233777 711197 233853 0 FreeSans 480 0 0 0 bidir_IE[21]
port 363 nsew
flabel metal3 710897 245234 711197 245310 0 FreeSans 480 0 0 0 bidir_SL[21]
port 409 nsew
flabel metal3 710897 245380 711197 245456 0 FreeSans 480 0 0 0 bidir_A[21]
port 455 nsew
flabel metal3 710897 245526 711197 245602 0 FreeSans 480 0 0 0 bidir_OE[21]
port 501 nsew
flabel metal3 710897 245672 711197 245748 0 FreeSans 480 0 0 0 bidir_Y[21]
port 547 nsew
flabel metal3 710897 247058 711197 247134 0 FreeSans 480 0 0 0 loopback_one[21]
port 599 nsew
flabel metal3 710897 247246 711197 247322 0 FreeSans 480 0 0 0 loopback_zero[21]
port 651 nsew
flabel metal3 710897 260372 711197 260448 0 FreeSans 480 0 0 0 bidir_CS[22]
port 86 nsew
flabel metal3 710897 260893 711197 260969 0 FreeSans 480 0 0 0 bidir_PU[22]
port 132 nsew
flabel metal3 710897 261122 711197 261198 0 FreeSans 480 0 0 0 bidir_PDRV0[22]
port 178 nsew
flabel metal3 710897 261264 711197 261340 0 FreeSans 480 0 0 0 bidir_PDRV1[22]
port 224 nsew
flabel metal3 710897 261406 711197 261482 0 FreeSans 480 0 0 0 bidir_ANA[22]
port 270 nsew
flabel metal3 710897 261766 711197 261842 0 FreeSans 480 0 0 0 bidir_PD[22]
port 316 nsew
flabel metal3 710897 261977 711197 262053 0 FreeSans 480 0 0 0 bidir_IE[22]
port 362 nsew
flabel metal3 710897 273434 711197 273510 0 FreeSans 480 0 0 0 bidir_SL[22]
port 408 nsew
flabel metal3 710897 273580 711197 273656 0 FreeSans 480 0 0 0 bidir_A[22]
port 454 nsew
flabel metal3 710897 273726 711197 273802 0 FreeSans 480 0 0 0 bidir_OE[22]
port 500 nsew
flabel metal3 710897 273872 711197 273948 0 FreeSans 480 0 0 0 bidir_Y[22]
port 546 nsew
flabel metal3 710897 275258 711197 275334 0 FreeSans 480 0 0 0 loopback_one[22]
port 598 nsew
flabel metal3 710897 275446 711197 275522 0 FreeSans 480 0 0 0 loopback_zero[22]
port 650 nsew
flabel metal3 710897 288572 711197 288648 0 FreeSans 480 0 0 0 bidir_CS[23]
port 85 nsew
flabel metal3 710897 289093 711197 289169 0 FreeSans 480 0 0 0 bidir_PU[23]
port 131 nsew
flabel metal3 710897 289322 711197 289398 0 FreeSans 480 0 0 0 bidir_PDRV0[23]
port 177 nsew
flabel metal3 710897 289464 711197 289540 0 FreeSans 480 0 0 0 bidir_PDRV1[23]
port 223 nsew
flabel metal3 710897 289606 711197 289682 0 FreeSans 480 0 0 0 bidir_ANA[23]
port 269 nsew
flabel metal3 710897 289966 711197 290042 0 FreeSans 480 0 0 0 bidir_PD[23]
port 315 nsew
flabel metal3 710897 290177 711197 290253 0 FreeSans 480 0 0 0 bidir_IE[23]
port 361 nsew
flabel metal3 710897 301634 711197 301710 0 FreeSans 480 0 0 0 bidir_SL[23]
port 407 nsew
flabel metal3 710897 301780 711197 301856 0 FreeSans 480 0 0 0 bidir_A[23]
port 453 nsew
flabel metal3 710897 301926 711197 302002 0 FreeSans 480 0 0 0 bidir_OE[23]
port 499 nsew
flabel metal3 710897 302072 711197 302148 0 FreeSans 480 0 0 0 bidir_Y[23]
port 545 nsew
flabel metal3 710897 303458 711197 303534 0 FreeSans 480 0 0 0 loopback_one[23]
port 597 nsew
flabel metal3 710897 303646 711197 303722 0 FreeSans 480 0 0 0 loopback_zero[23]
port 649 nsew
flabel metal3 710897 316772 711197 316848 0 FreeSans 480 0 0 0 bidir_CS[24]
port 84 nsew
flabel metal3 710897 317293 711197 317369 0 FreeSans 480 0 0 0 bidir_PU[24]
port 130 nsew
flabel metal3 710897 317522 711197 317598 0 FreeSans 480 0 0 0 bidir_PDRV0[24]
port 176 nsew
flabel metal3 710897 317664 711197 317740 0 FreeSans 480 0 0 0 bidir_PDRV1[24]
port 222 nsew
flabel metal3 710897 317806 711197 317882 0 FreeSans 480 0 0 0 bidir_ANA[24]
port 268 nsew
flabel metal3 710897 318166 711197 318242 0 FreeSans 480 0 0 0 bidir_PD[24]
port 314 nsew
flabel metal3 710897 318377 711197 318453 0 FreeSans 480 0 0 0 bidir_IE[24]
port 360 nsew
flabel metal3 710897 329834 711197 329910 0 FreeSans 480 0 0 0 bidir_SL[24]
port 406 nsew
flabel metal3 710897 329980 711197 330056 0 FreeSans 480 0 0 0 bidir_A[24]
port 452 nsew
flabel metal3 710897 330126 711197 330202 0 FreeSans 480 0 0 0 bidir_OE[24]
port 498 nsew
flabel metal3 710897 330272 711197 330348 0 FreeSans 480 0 0 0 bidir_Y[24]
port 544 nsew
flabel metal3 710897 331658 711197 331734 0 FreeSans 480 0 0 0 loopback_one[24]
port 596 nsew
flabel metal3 710897 331846 711197 331922 0 FreeSans 480 0 0 0 loopback_zero[24]
port 648 nsew
flabel metal3 710897 344972 711197 345048 0 FreeSans 480 0 0 0 bidir_CS[25]
port 83 nsew
flabel metal3 710897 345493 711197 345569 0 FreeSans 480 0 0 0 bidir_PU[25]
port 129 nsew
flabel metal3 710897 345722 711197 345798 0 FreeSans 480 0 0 0 bidir_PDRV0[25]
port 175 nsew
flabel metal3 710897 345864 711197 345940 0 FreeSans 480 0 0 0 bidir_PDRV1[25]
port 221 nsew
flabel metal3 710897 346006 711197 346082 0 FreeSans 480 0 0 0 bidir_ANA[25]
port 267 nsew
flabel metal3 710897 346366 711197 346442 0 FreeSans 480 0 0 0 bidir_PD[25]
port 313 nsew
flabel metal3 710897 346577 711197 346653 0 FreeSans 480 0 0 0 bidir_IE[25]
port 359 nsew
flabel metal3 710897 358034 711197 358110 0 FreeSans 480 0 0 0 bidir_SL[25]
port 405 nsew
flabel metal3 710897 358180 711197 358256 0 FreeSans 480 0 0 0 bidir_A[25]
port 451 nsew
flabel metal3 710897 358326 711197 358402 0 FreeSans 480 0 0 0 bidir_OE[25]
port 497 nsew
flabel metal3 710897 358472 711197 358548 0 FreeSans 480 0 0 0 bidir_Y[25]
port 543 nsew
flabel metal3 710897 359858 711197 359934 0 FreeSans 480 0 0 0 loopback_one[25]
port 595 nsew
flabel metal3 710897 360046 711197 360122 0 FreeSans 480 0 0 0 loopback_zero[25]
port 647 nsew
flabel metal2 683072 430768 683148 431068 0 FreeSans 480 90 0 0 bidir_CS[26]
port 82 nsew
flabel metal2 683593 430768 683669 431068 0 FreeSans 480 90 0 0 bidir_PU[26]
port 128 nsew
flabel metal2 683822 430768 683898 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[26]
port 174 nsew
flabel metal2 683964 430768 684040 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[26]
port 220 nsew
flabel metal2 684106 430768 684182 431068 0 FreeSans 480 90 0 0 bidir_ANA[26]
port 266 nsew
flabel metal2 684466 430768 684542 431068 0 FreeSans 480 90 0 0 bidir_PD[26]
port 312 nsew
flabel metal2 684677 430768 684753 431068 0 FreeSans 480 90 0 0 bidir_IE[26]
port 358 nsew
flabel metal2 696134 430768 696210 431068 0 FreeSans 480 90 0 0 bidir_SL[26]
port 404 nsew
flabel metal2 696280 430768 696356 431068 0 FreeSans 480 90 0 0 bidir_A[26]
port 450 nsew
flabel metal2 696426 430768 696502 431068 0 FreeSans 480 90 0 0 bidir_OE[26]
port 496 nsew
flabel metal2 696572 430768 696648 431068 0 FreeSans 480 90 0 0 bidir_Y[26]
port 542 nsew
flabel metal2 697958 430768 698034 431068 0 FreeSans 480 90 0 0 loopback_one[26]
port 594 nsew
flabel metal2 698146 430768 698222 431068 0 FreeSans 480 90 0 0 loopback_zero[26]
port 646 nsew
flabel metal2 657272 430768 657348 431068 0 FreeSans 480 90 0 0 bidir_CS[27]
port 81 nsew
flabel metal2 657793 430768 657869 431068 0 FreeSans 480 90 0 0 bidir_PU[27]
port 127 nsew
flabel metal2 658022 430768 658098 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[27]
port 173 nsew
flabel metal2 658164 430768 658240 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[27]
port 219 nsew
flabel metal2 658306 430768 658382 431068 0 FreeSans 480 90 0 0 bidir_ANA[27]
port 265 nsew
flabel metal2 658666 430768 658742 431068 0 FreeSans 480 90 0 0 bidir_PD[27]
port 311 nsew
flabel metal2 658877 430768 658953 431068 0 FreeSans 480 90 0 0 bidir_IE[27]
port 357 nsew
flabel metal2 670334 430768 670410 431068 0 FreeSans 480 90 0 0 bidir_SL[27]
port 403 nsew
flabel metal2 670480 430768 670556 431068 0 FreeSans 480 90 0 0 bidir_A[27]
port 449 nsew
flabel metal2 670626 430768 670702 431068 0 FreeSans 480 90 0 0 bidir_OE[27]
port 495 nsew
flabel metal2 670772 430768 670848 431068 0 FreeSans 480 90 0 0 bidir_Y[27]
port 541 nsew
flabel metal2 672158 430768 672234 431068 0 FreeSans 480 90 0 0 loopback_one[27]
port 593 nsew
flabel metal2 672346 430768 672422 431068 0 FreeSans 480 90 0 0 loopback_zero[27]
port 645 nsew
flabel metal2 631472 430768 631548 431068 0 FreeSans 480 90 0 0 bidir_CS[28]
port 80 nsew
flabel metal2 631993 430768 632069 431068 0 FreeSans 480 90 0 0 bidir_PU[28]
port 126 nsew
flabel metal2 632222 430768 632298 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[28]
port 172 nsew
flabel metal2 632364 430768 632440 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[28]
port 218 nsew
flabel metal2 632506 430768 632582 431068 0 FreeSans 480 90 0 0 bidir_ANA[28]
port 264 nsew
flabel metal2 632866 430768 632942 431068 0 FreeSans 480 90 0 0 bidir_PD[28]
port 310 nsew
flabel metal2 633077 430768 633153 431068 0 FreeSans 480 90 0 0 bidir_IE[28]
port 356 nsew
flabel metal2 644534 430768 644610 431068 0 FreeSans 480 90 0 0 bidir_SL[28]
port 402 nsew
flabel metal2 644680 430768 644756 431068 0 FreeSans 480 90 0 0 bidir_A[28]
port 448 nsew
flabel metal2 644826 430768 644902 431068 0 FreeSans 480 90 0 0 bidir_OE[28]
port 494 nsew
flabel metal2 644972 430768 645048 431068 0 FreeSans 480 90 0 0 bidir_Y[28]
port 540 nsew
flabel metal2 646358 430768 646434 431068 0 FreeSans 480 90 0 0 loopback_one[28]
port 592 nsew
flabel metal2 646546 430768 646622 431068 0 FreeSans 480 90 0 0 loopback_zero[28]
port 644 nsew
flabel metal2 605672 430768 605748 431068 0 FreeSans 480 90 0 0 bidir_CS[29]
port 79 nsew
flabel metal2 606193 430768 606269 431068 0 FreeSans 480 90 0 0 bidir_PU[29]
port 125 nsew
flabel metal2 606422 430768 606498 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[29]
port 171 nsew
flabel metal2 606564 430768 606640 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[29]
port 217 nsew
flabel metal2 606706 430768 606782 431068 0 FreeSans 480 90 0 0 bidir_ANA[29]
port 263 nsew
flabel metal2 607066 430768 607142 431068 0 FreeSans 480 90 0 0 bidir_PD[29]
port 309 nsew
flabel metal2 607277 430768 607353 431068 0 FreeSans 480 90 0 0 bidir_IE[29]
port 355 nsew
flabel metal2 618734 430768 618810 431068 0 FreeSans 480 90 0 0 bidir_SL[29]
port 401 nsew
flabel metal2 618880 430768 618956 431068 0 FreeSans 480 90 0 0 bidir_A[29]
port 447 nsew
flabel metal2 619026 430768 619102 431068 0 FreeSans 480 90 0 0 bidir_OE[29]
port 493 nsew
flabel metal2 619172 430768 619248 431068 0 FreeSans 480 90 0 0 bidir_Y[29]
port 539 nsew
flabel metal2 620558 430768 620634 431068 0 FreeSans 480 90 0 0 loopback_one[29]
port 591 nsew
flabel metal2 620746 430768 620822 431068 0 FreeSans 480 90 0 0 loopback_zero[29]
port 643 nsew
flabel metal2 528272 430768 528348 431068 0 FreeSans 480 90 0 0 bidir_CS[30]
port 78 nsew
flabel metal2 528793 430768 528869 431068 0 FreeSans 480 90 0 0 bidir_PU[30]
port 124 nsew
flabel metal2 529022 430768 529098 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[30]
port 170 nsew
flabel metal2 529164 430768 529240 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[30]
port 216 nsew
flabel metal2 529306 430768 529382 431068 0 FreeSans 480 90 0 0 bidir_ANA[30]
port 262 nsew
flabel metal2 529666 430768 529742 431068 0 FreeSans 480 90 0 0 bidir_PD[30]
port 308 nsew
flabel metal2 529877 430768 529953 431068 0 FreeSans 480 90 0 0 bidir_IE[30]
port 354 nsew
flabel metal2 541334 430768 541410 431068 0 FreeSans 480 90 0 0 bidir_SL[30]
port 400 nsew
flabel metal2 541480 430768 541556 431068 0 FreeSans 480 90 0 0 bidir_A[30]
port 446 nsew
flabel metal2 541626 430768 541702 431068 0 FreeSans 480 90 0 0 bidir_OE[30]
port 492 nsew
flabel metal2 541772 430768 541848 431068 0 FreeSans 480 90 0 0 bidir_Y[30]
port 538 nsew
flabel metal2 543158 430768 543234 431068 0 FreeSans 480 90 0 0 loopback_one[30]
port 590 nsew
flabel metal2 543346 430768 543422 431068 0 FreeSans 480 90 0 0 loopback_zero[30]
port 642 nsew
flabel metal2 502472 430768 502548 431068 0 FreeSans 480 90 0 0 bidir_CS[31]
port 77 nsew
flabel metal2 502993 430768 503069 431068 0 FreeSans 480 90 0 0 bidir_PU[31]
port 123 nsew
flabel metal2 503222 430768 503298 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[31]
port 169 nsew
flabel metal2 503364 430768 503440 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[31]
port 215 nsew
flabel metal2 503506 430768 503582 431068 0 FreeSans 480 90 0 0 bidir_ANA[31]
port 261 nsew
flabel metal2 503866 430768 503942 431068 0 FreeSans 480 90 0 0 bidir_PD[31]
port 307 nsew
flabel metal2 504077 430768 504153 431068 0 FreeSans 480 90 0 0 bidir_IE[31]
port 353 nsew
flabel metal2 515534 430768 515610 431068 0 FreeSans 480 90 0 0 bidir_SL[31]
port 399 nsew
flabel metal2 515680 430768 515756 431068 0 FreeSans 480 90 0 0 bidir_A[31]
port 445 nsew
flabel metal2 515826 430768 515902 431068 0 FreeSans 480 90 0 0 bidir_OE[31]
port 491 nsew
flabel metal2 515972 430768 516048 431068 0 FreeSans 480 90 0 0 bidir_Y[31]
port 537 nsew
flabel metal2 517358 430768 517434 431068 0 FreeSans 480 90 0 0 loopback_one[31]
port 589 nsew
flabel metal2 517546 430768 517622 431068 0 FreeSans 480 90 0 0 loopback_zero[31]
port 641 nsew
flabel metal2 476672 430768 476748 431068 0 FreeSans 480 90 0 0 bidir_CS[32]
port 76 nsew
flabel metal2 477193 430768 477269 431068 0 FreeSans 480 90 0 0 bidir_PU[32]
port 122 nsew
flabel metal2 477422 430768 477498 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[32]
port 168 nsew
flabel metal2 477564 430768 477640 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[32]
port 214 nsew
flabel metal2 477706 430768 477782 431068 0 FreeSans 480 90 0 0 bidir_ANA[32]
port 260 nsew
flabel metal2 478066 430768 478142 431068 0 FreeSans 480 90 0 0 bidir_PD[32]
port 306 nsew
flabel metal2 478277 430768 478353 431068 0 FreeSans 480 90 0 0 bidir_IE[32]
port 352 nsew
flabel metal2 489734 430768 489810 431068 0 FreeSans 480 90 0 0 bidir_SL[32]
port 398 nsew
flabel metal2 489880 430768 489956 431068 0 FreeSans 480 90 0 0 bidir_A[32]
port 444 nsew
flabel metal2 490026 430768 490102 431068 0 FreeSans 480 90 0 0 bidir_OE[32]
port 490 nsew
flabel metal2 490172 430768 490248 431068 0 FreeSans 480 90 0 0 bidir_Y[32]
port 536 nsew
flabel metal2 491558 430768 491634 431068 0 FreeSans 480 90 0 0 loopback_one[32]
port 588 nsew
flabel metal2 491746 430768 491822 431068 0 FreeSans 480 90 0 0 loopback_zero[32]
port 640 nsew
flabel metal2 450872 430768 450948 431068 0 FreeSans 480 90 0 0 bidir_CS[33]
port 75 nsew
flabel metal2 451393 430768 451469 431068 0 FreeSans 480 90 0 0 bidir_PU[33]
port 121 nsew
flabel metal2 451622 430768 451698 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[33]
port 167 nsew
flabel metal2 451764 430768 451840 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[33]
port 213 nsew
flabel metal2 451906 430768 451982 431068 0 FreeSans 480 90 0 0 bidir_ANA[33]
port 259 nsew
flabel metal2 452266 430768 452342 431068 0 FreeSans 480 90 0 0 bidir_PD[33]
port 305 nsew
flabel metal2 452477 430768 452553 431068 0 FreeSans 480 90 0 0 bidir_IE[33]
port 351 nsew
flabel metal2 463934 430768 464010 431068 0 FreeSans 480 90 0 0 bidir_SL[33]
port 397 nsew
flabel metal2 464080 430768 464156 431068 0 FreeSans 480 90 0 0 bidir_A[33]
port 443 nsew
flabel metal2 464226 430768 464302 431068 0 FreeSans 480 90 0 0 bidir_OE[33]
port 489 nsew
flabel metal2 464372 430768 464448 431068 0 FreeSans 480 90 0 0 bidir_Y[33]
port 535 nsew
flabel metal2 465758 430768 465834 431068 0 FreeSans 480 90 0 0 loopback_one[33]
port 587 nsew
flabel metal2 465946 430768 466022 431068 0 FreeSans 480 90 0 0 loopback_zero[33]
port 639 nsew
flabel metal2 425072 430768 425148 431068 0 FreeSans 480 90 0 0 bidir_CS[34]
port 74 nsew
flabel metal2 425593 430768 425669 431068 0 FreeSans 480 90 0 0 bidir_PU[34]
port 120 nsew
flabel metal2 425822 430768 425898 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[34]
port 166 nsew
flabel metal2 425964 430768 426040 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[34]
port 212 nsew
flabel metal2 426106 430768 426182 431068 0 FreeSans 480 90 0 0 bidir_ANA[34]
port 258 nsew
flabel metal2 426466 430768 426542 431068 0 FreeSans 480 90 0 0 bidir_PD[34]
port 304 nsew
flabel metal2 426677 430768 426753 431068 0 FreeSans 480 90 0 0 bidir_IE[34]
port 350 nsew
flabel metal2 438134 430768 438210 431068 0 FreeSans 480 90 0 0 bidir_SL[34]
port 396 nsew
flabel metal2 438280 430768 438356 431068 0 FreeSans 480 90 0 0 bidir_A[34]
port 442 nsew
flabel metal2 438426 430768 438502 431068 0 FreeSans 480 90 0 0 bidir_OE[34]
port 488 nsew
flabel metal2 438572 430768 438648 431068 0 FreeSans 480 90 0 0 bidir_Y[34]
port 534 nsew
flabel metal2 439958 430768 440034 431068 0 FreeSans 480 90 0 0 loopback_one[34]
port 586 nsew
flabel metal2 440146 430768 440222 431068 0 FreeSans 480 90 0 0 loopback_zero[34]
port 638 nsew
flabel metal2 399272 430768 399348 431068 0 FreeSans 480 90 0 0 bidir_CS[35]
port 73 nsew
flabel metal2 399793 430768 399869 431068 0 FreeSans 480 90 0 0 bidir_PU[35]
port 119 nsew
flabel metal2 400022 430768 400098 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[35]
port 165 nsew
flabel metal2 400164 430768 400240 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[35]
port 211 nsew
flabel metal2 400306 430768 400382 431068 0 FreeSans 480 90 0 0 bidir_ANA[35]
port 257 nsew
flabel metal2 400666 430768 400742 431068 0 FreeSans 480 90 0 0 bidir_PD[35]
port 303 nsew
flabel metal2 400877 430768 400953 431068 0 FreeSans 480 90 0 0 bidir_IE[35]
port 349 nsew
flabel metal2 412334 430768 412410 431068 0 FreeSans 480 90 0 0 bidir_SL[35]
port 395 nsew
flabel metal2 412480 430768 412556 431068 0 FreeSans 480 90 0 0 bidir_A[35]
port 441 nsew
flabel metal2 412626 430768 412702 431068 0 FreeSans 480 90 0 0 bidir_OE[35]
port 487 nsew
flabel metal2 412772 430768 412848 431068 0 FreeSans 480 90 0 0 bidir_Y[35]
port 533 nsew
flabel metal2 414158 430768 414234 431068 0 FreeSans 480 90 0 0 loopback_one[35]
port 585 nsew
flabel metal2 414346 430768 414422 431068 0 FreeSans 480 90 0 0 loopback_zero[35]
port 637 nsew
flabel metal2 373472 430768 373548 431068 0 FreeSans 480 90 0 0 bidir_CS[36]
port 72 nsew
flabel metal2 373993 430768 374069 431068 0 FreeSans 480 90 0 0 bidir_PU[36]
port 118 nsew
flabel metal2 374222 430768 374298 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[36]
port 164 nsew
flabel metal2 374364 430768 374440 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[36]
port 210 nsew
flabel metal2 374506 430768 374582 431068 0 FreeSans 480 90 0 0 bidir_ANA[36]
port 256 nsew
flabel metal2 374866 430768 374942 431068 0 FreeSans 480 90 0 0 bidir_PD[36]
port 302 nsew
flabel metal2 375077 430768 375153 431068 0 FreeSans 480 90 0 0 bidir_IE[36]
port 348 nsew
flabel metal2 386534 430768 386610 431068 0 FreeSans 480 90 0 0 bidir_SL[36]
port 394 nsew
flabel metal2 386680 430768 386756 431068 0 FreeSans 480 90 0 0 bidir_A[36]
port 440 nsew
flabel metal2 386826 430768 386902 431068 0 FreeSans 480 90 0 0 bidir_OE[36]
port 486 nsew
flabel metal2 386972 430768 387048 431068 0 FreeSans 480 90 0 0 bidir_Y[36]
port 532 nsew
flabel metal2 388358 430768 388434 431068 0 FreeSans 480 90 0 0 loopback_one[36]
port 584 nsew
flabel metal2 388546 430768 388622 431068 0 FreeSans 480 90 0 0 loopback_zero[36]
port 636 nsew
flabel metal2 347672 430768 347748 431068 0 FreeSans 480 90 0 0 bidir_CS[37]
port 71 nsew
flabel metal2 348193 430768 348269 431068 0 FreeSans 480 90 0 0 bidir_PU[37]
port 117 nsew
flabel metal2 348422 430768 348498 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[37]
port 163 nsew
flabel metal2 348564 430768 348640 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[37]
port 209 nsew
flabel metal2 348706 430768 348782 431068 0 FreeSans 480 90 0 0 bidir_ANA[37]
port 255 nsew
flabel metal2 349066 430768 349142 431068 0 FreeSans 480 90 0 0 bidir_PD[37]
port 301 nsew
flabel metal2 349277 430768 349353 431068 0 FreeSans 480 90 0 0 bidir_IE[37]
port 347 nsew
flabel metal2 360734 430768 360810 431068 0 FreeSans 480 90 0 0 bidir_SL[37]
port 393 nsew
flabel metal2 360880 430768 360956 431068 0 FreeSans 480 90 0 0 bidir_A[37]
port 439 nsew
flabel metal2 361026 430768 361102 431068 0 FreeSans 480 90 0 0 bidir_OE[37]
port 485 nsew
flabel metal2 361172 430768 361248 431068 0 FreeSans 480 90 0 0 bidir_Y[37]
port 531 nsew
flabel metal2 362558 430768 362634 431068 0 FreeSans 480 90 0 0 loopback_one[37]
port 583 nsew
flabel metal2 362746 430768 362822 431068 0 FreeSans 480 90 0 0 loopback_zero[37]
port 635 nsew
flabel metal2 321872 430768 321948 431068 0 FreeSans 480 90 0 0 bidir_CS[38]
port 70 nsew
flabel metal2 322393 430768 322469 431068 0 FreeSans 480 90 0 0 bidir_PU[38]
port 116 nsew
flabel metal2 322622 430768 322698 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[38]
port 162 nsew
flabel metal2 322764 430768 322840 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[38]
port 208 nsew
flabel metal2 322906 430768 322982 431068 0 FreeSans 480 90 0 0 bidir_ANA[38]
port 254 nsew
flabel metal2 323266 430768 323342 431068 0 FreeSans 480 90 0 0 bidir_PD[38]
port 300 nsew
flabel metal2 323477 430768 323553 431068 0 FreeSans 480 90 0 0 bidir_IE[38]
port 346 nsew
flabel metal2 334934 430768 335010 431068 0 FreeSans 480 90 0 0 bidir_SL[38]
port 392 nsew
flabel metal2 335080 430768 335156 431068 0 FreeSans 480 90 0 0 bidir_A[38]
port 438 nsew
flabel metal2 335226 430768 335302 431068 0 FreeSans 480 90 0 0 bidir_OE[38]
port 484 nsew
flabel metal2 335372 430768 335448 431068 0 FreeSans 480 90 0 0 bidir_Y[38]
port 530 nsew
flabel metal2 336758 430768 336834 431068 0 FreeSans 480 90 0 0 loopback_one[38]
port 582 nsew
flabel metal2 336946 430768 337022 431068 0 FreeSans 480 90 0 0 loopback_zero[38]
port 634 nsew
flabel metal2 296072 430768 296148 431068 0 FreeSans 480 90 0 0 bidir_CS[39]
port 69 nsew
flabel metal2 296593 430768 296669 431068 0 FreeSans 480 90 0 0 bidir_PU[39]
port 115 nsew
flabel metal2 296822 430768 296898 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[39]
port 161 nsew
flabel metal2 296964 430768 297040 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[39]
port 207 nsew
flabel metal2 297106 430768 297182 431068 0 FreeSans 480 90 0 0 bidir_ANA[39]
port 253 nsew
flabel metal2 297466 430768 297542 431068 0 FreeSans 480 90 0 0 bidir_PD[39]
port 299 nsew
flabel metal2 297677 430768 297753 431068 0 FreeSans 480 90 0 0 bidir_IE[39]
port 345 nsew
flabel metal2 309134 430768 309210 431068 0 FreeSans 480 90 0 0 bidir_SL[39]
port 391 nsew
flabel metal2 309280 430768 309356 431068 0 FreeSans 480 90 0 0 bidir_A[39]
port 437 nsew
flabel metal2 309426 430768 309502 431068 0 FreeSans 480 90 0 0 bidir_OE[39]
port 483 nsew
flabel metal2 309572 430768 309648 431068 0 FreeSans 480 90 0 0 bidir_Y[39]
port 529 nsew
flabel metal2 310958 430768 311034 431068 0 FreeSans 480 90 0 0 loopback_one[39]
port 581 nsew
flabel metal2 311146 430768 311222 431068 0 FreeSans 480 90 0 0 loopback_zero[39]
port 633 nsew
flabel metal2 270272 430768 270348 431068 0 FreeSans 480 90 0 0 bidir_CS[40]
port 68 nsew
flabel metal2 270793 430768 270869 431068 0 FreeSans 480 90 0 0 bidir_PU[40]
port 114 nsew
flabel metal2 271022 430768 271098 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[40]
port 160 nsew
flabel metal2 271164 430768 271240 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[40]
port 206 nsew
flabel metal2 271306 430768 271382 431068 0 FreeSans 480 90 0 0 bidir_ANA[40]
port 252 nsew
flabel metal2 271666 430768 271742 431068 0 FreeSans 480 90 0 0 bidir_PD[40]
port 298 nsew
flabel metal2 271877 430768 271953 431068 0 FreeSans 480 90 0 0 bidir_IE[40]
port 344 nsew
flabel metal2 283334 430768 283410 431068 0 FreeSans 480 90 0 0 bidir_SL[40]
port 390 nsew
flabel metal2 283480 430768 283556 431068 0 FreeSans 480 90 0 0 bidir_A[40]
port 436 nsew
flabel metal2 283626 430768 283702 431068 0 FreeSans 480 90 0 0 bidir_OE[40]
port 482 nsew
flabel metal2 283772 430768 283848 431068 0 FreeSans 480 90 0 0 bidir_Y[40]
port 528 nsew
flabel metal2 285158 430768 285234 431068 0 FreeSans 480 90 0 0 loopback_one[40]
port 580 nsew
flabel metal2 285346 430768 285422 431068 0 FreeSans 480 90 0 0 loopback_zero[40]
port 632 nsew
flabel metal2 244472 430768 244548 431068 0 FreeSans 480 90 0 0 bidir_CS[41]
port 67 nsew
flabel metal2 244993 430768 245069 431068 0 FreeSans 480 90 0 0 bidir_PU[41]
port 113 nsew
flabel metal2 245222 430768 245298 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[41]
port 159 nsew
flabel metal2 245364 430768 245440 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[41]
port 205 nsew
flabel metal2 245506 430768 245582 431068 0 FreeSans 480 90 0 0 bidir_ANA[41]
port 251 nsew
flabel metal2 245866 430768 245942 431068 0 FreeSans 480 90 0 0 bidir_PD[41]
port 297 nsew
flabel metal2 246077 430768 246153 431068 0 FreeSans 480 90 0 0 bidir_IE[41]
port 343 nsew
flabel metal2 257534 430768 257610 431068 0 FreeSans 480 90 0 0 bidir_SL[41]
port 389 nsew
flabel metal2 257680 430768 257756 431068 0 FreeSans 480 90 0 0 bidir_A[41]
port 435 nsew
flabel metal2 257826 430768 257902 431068 0 FreeSans 480 90 0 0 bidir_OE[41]
port 481 nsew
flabel metal2 257972 430768 258048 431068 0 FreeSans 480 90 0 0 bidir_Y[41]
port 527 nsew
flabel metal2 259358 430768 259434 431068 0 FreeSans 480 90 0 0 loopback_one[41]
port 579 nsew
flabel metal2 259546 430768 259622 431068 0 FreeSans 480 90 0 0 loopback_zero[41]
port 631 nsew
flabel metal2 167072 430768 167148 431068 0 FreeSans 480 90 0 0 bidir_CS[42]
port 66 nsew
flabel metal2 167593 430768 167669 431068 0 FreeSans 480 90 0 0 bidir_PU[42]
port 112 nsew
flabel metal2 167822 430768 167898 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[42]
port 158 nsew
flabel metal2 167964 430768 168040 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[42]
port 204 nsew
flabel metal2 168106 430768 168182 431068 0 FreeSans 480 90 0 0 bidir_ANA[42]
port 250 nsew
flabel metal2 168466 430768 168542 431068 0 FreeSans 480 90 0 0 bidir_PD[42]
port 296 nsew
flabel metal2 168677 430768 168753 431068 0 FreeSans 480 90 0 0 bidir_IE[42]
port 342 nsew
flabel metal2 180134 430768 180210 431068 0 FreeSans 480 90 0 0 bidir_SL[42]
port 388 nsew
flabel metal2 180280 430768 180356 431068 0 FreeSans 480 90 0 0 bidir_A[42]
port 434 nsew
flabel metal2 180426 430768 180502 431068 0 FreeSans 480 90 0 0 bidir_OE[42]
port 480 nsew
flabel metal2 180572 430768 180648 431068 0 FreeSans 480 90 0 0 bidir_Y[42]
port 526 nsew
flabel metal2 181958 430768 182034 431068 0 FreeSans 480 90 0 0 loopback_one[42]
port 578 nsew
flabel metal2 182146 430768 182222 431068 0 FreeSans 480 90 0 0 loopback_zero[42]
port 630 nsew
flabel metal2 141272 430768 141348 431068 0 FreeSans 480 90 0 0 bidir_CS[43]
port 65 nsew
flabel metal2 141793 430768 141869 431068 0 FreeSans 480 90 0 0 bidir_PU[43]
port 111 nsew
flabel metal2 142022 430768 142098 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[43]
port 157 nsew
flabel metal2 142164 430768 142240 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[43]
port 203 nsew
flabel metal2 142306 430768 142382 431068 0 FreeSans 480 90 0 0 bidir_ANA[43]
port 249 nsew
flabel metal2 142666 430768 142742 431068 0 FreeSans 480 90 0 0 bidir_PD[43]
port 295 nsew
flabel metal2 142877 430768 142953 431068 0 FreeSans 480 90 0 0 bidir_IE[43]
port 341 nsew
flabel metal2 154334 430768 154410 431068 0 FreeSans 480 90 0 0 bidir_SL[43]
port 387 nsew
flabel metal2 154480 430768 154556 431068 0 FreeSans 480 90 0 0 bidir_A[43]
port 433 nsew
flabel metal2 154626 430768 154702 431068 0 FreeSans 480 90 0 0 bidir_OE[43]
port 479 nsew
flabel metal2 154772 430768 154848 431068 0 FreeSans 480 90 0 0 bidir_Y[43]
port 525 nsew
flabel metal2 156158 430768 156234 431068 0 FreeSans 480 90 0 0 loopback_one[43]
port 577 nsew
flabel metal2 156346 430768 156422 431068 0 FreeSans 480 90 0 0 loopback_zero[43]
port 629 nsew
flabel metal2 115472 430768 115548 431068 0 FreeSans 480 90 0 0 bidir_CS[44]
port 64 nsew
flabel metal2 115993 430768 116069 431068 0 FreeSans 480 90 0 0 bidir_PU[44]
port 110 nsew
flabel metal2 116222 430768 116298 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[44]
port 156 nsew
flabel metal2 116364 430768 116440 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[44]
port 202 nsew
flabel metal2 116506 430768 116582 431068 0 FreeSans 480 90 0 0 bidir_ANA[44]
port 248 nsew
flabel metal2 116866 430768 116942 431068 0 FreeSans 480 90 0 0 bidir_PD[44]
port 294 nsew
flabel metal2 117077 430768 117153 431068 0 FreeSans 480 90 0 0 bidir_IE[44]
port 340 nsew
flabel metal2 128534 430768 128610 431068 0 FreeSans 480 90 0 0 bidir_SL[44]
port 386 nsew
flabel metal2 128680 430768 128756 431068 0 FreeSans 480 90 0 0 bidir_A[44]
port 432 nsew
flabel metal2 128826 430768 128902 431068 0 FreeSans 480 90 0 0 bidir_OE[44]
port 478 nsew
flabel metal2 128972 430768 129048 431068 0 FreeSans 480 90 0 0 bidir_Y[44]
port 524 nsew
flabel metal2 130358 430768 130434 431068 0 FreeSans 480 90 0 0 loopback_one[44]
port 576 nsew
flabel metal2 130546 430768 130622 431068 0 FreeSans 480 90 0 0 loopback_zero[44]
port 628 nsew
flabel metal2 89672 430768 89748 431068 0 FreeSans 480 90 0 0 bidir_CS[45]
port 63 nsew
flabel metal2 90193 430768 90269 431068 0 FreeSans 480 90 0 0 bidir_PU[45]
port 109 nsew
flabel metal2 90422 430768 90498 431068 0 FreeSans 480 90 0 0 bidir_PDRV0[45]
port 155 nsew
flabel metal2 90564 430768 90640 431068 0 FreeSans 480 90 0 0 bidir_PDRV1[45]
port 201 nsew
flabel metal2 90706 430768 90782 431068 0 FreeSans 480 90 0 0 bidir_ANA[45]
port 247 nsew
flabel metal2 91066 430768 91142 431068 0 FreeSans 480 90 0 0 bidir_PD[45]
port 293 nsew
flabel metal2 91277 430768 91353 431068 0 FreeSans 480 90 0 0 bidir_IE[45]
port 339 nsew
flabel metal2 102734 430768 102810 431068 0 FreeSans 480 90 0 0 bidir_SL[45]
port 385 nsew
flabel metal2 102880 430768 102956 431068 0 FreeSans 480 90 0 0 bidir_A[45]
port 431 nsew
flabel metal2 103026 430768 103102 431068 0 FreeSans 480 90 0 0 bidir_OE[45]
port 477 nsew
flabel metal2 103172 430768 103248 431068 0 FreeSans 480 90 0 0 bidir_Y[45]
port 523 nsew
flabel metal2 104558 430768 104634 431068 0 FreeSans 480 90 0 0 loopback_one[45]
port 575 nsew
flabel metal2 104746 430768 104822 431068 0 FreeSans 480 90 0 0 loopback_zero[45]
port 627 nsew
flabel metal3 75203 216158 75503 216234 0 FreeSans 480 0 0 0 input_PD[1]
port 681 nsew
flabel metal3 75203 217031 75503 217107 0 FreeSans 480 0 0 0 input_PU[1]
port 676 nsew
flabel metal3 75203 204052 75503 204128 0 FreeSans 480 0 0 0 input_Y[1]
port 686 nsew
flabel metal3 75203 232252 75503 232328 0 FreeSans 480 0 0 0 input_Y[0]
port 687 nsew
flabel metal3 75203 245231 75503 245307 0 FreeSans 480 0 0 0 input_PU[0]
port 677 nsew
flabel metal3 75203 244358 75503 244434 0 FreeSans 480 0 0 0 input_PD[0]
port 682 nsew
flabel metal3 75203 188831 75503 188907 0 FreeSans 480 0 0 0 input_PU[2]
port 675 nsew
flabel metal3 75203 187958 75503 188034 0 FreeSans 480 0 0 0 input_PD[2]
port 680 nsew
flabel metal3 75203 175852 75503 175928 0 FreeSans 480 0 0 0 input_Y[2]
port 685 nsew
flabel metal3 75203 160631 75503 160707 0 FreeSans 480 0 0 0 input_PU[3]
port 674 nsew
flabel metal3 75203 159758 75503 159834 0 FreeSans 480 0 0 0 input_PD[3]
port 679 nsew
flabel metal3 75203 147652 75503 147728 0 FreeSans 480 0 0 0 input_Y[3]
port 684 nsew
flabel metal3 75203 162458 75503 162534 0 FreeSans 480 0 0 0 loopback_one[49]
port 571 nsew
flabel metal3 75203 162646 75503 162722 0 FreeSans 480 0 0 0 loopback_zero[49]
port 623 nsew
flabel metal3 75203 190846 75503 190922 0 FreeSans 480 0 0 0 loopback_zero[48]
port 624 nsew
flabel metal3 75203 190658 75503 190734 0 FreeSans 480 0 0 0 loopback_one[48]
port 572 nsew
flabel metal3 75203 218858 75503 218934 0 FreeSans 480 0 0 0 loopback_one[47]
port 573 nsew
flabel metal3 75203 219046 75503 219122 0 FreeSans 480 0 0 0 loopback_zero[47]
port 625 nsew
flabel metal3 75203 247246 75503 247322 0 FreeSans 480 0 0 0 loopback_zero[46]
port 626 nsew
flabel metal3 75203 247058 75503 247134 0 FreeSans 480 0 0 0 loopback_one[46]
port 574 nsew
flabel metal2 74951 355724 75251 356232 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 354588 75251 355096 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 353452 75251 353960 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 352316 75251 352824 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 350776 75251 351284 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 349640 75251 350148 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 348504 75251 349012 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 347368 75251 347876 0 FreeSans 480 0 0 0 analog_PAD[0]
port 55 nsew
flabel metal2 74951 327524 75251 328032 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 326388 75251 326896 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 325252 75251 325760 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 324116 75251 324624 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 322576 75251 323084 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 321440 75251 321948 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 320304 75251 320812 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 319168 75251 319676 0 FreeSans 480 0 0 0 analog_PAD[1]
port 54 nsew
flabel metal2 74951 299324 75251 299832 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 298188 75251 298696 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 297052 75251 297560 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 295916 75251 296424 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 294376 75251 294884 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 293240 75251 293748 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 292104 75251 292612 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 290968 75251 291476 0 FreeSans 480 0 0 0 analog_PAD[2]
port 53 nsew
flabel metal2 74951 271124 75251 271632 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 269988 75251 270496 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 268852 75251 269360 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 267716 75251 268224 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 266176 75251 266684 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 265040 75251 265548 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 263904 75251 264412 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal2 74951 262768 75251 263276 0 FreeSans 480 0 0 0 analog_PAD[3]
port 52 nsew
flabel metal4 192474 75200 194370 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 194954 75200 197000 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 197324 75200 199370 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 200030 75200 202076 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 202400 75200 204446 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 205030 75200 206926 75400 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 218274 75200 220170 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 220754 75200 222800 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 223124 75200 225170 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 225830 75200 227876 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 228200 75200 230246 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 230830 75200 232726 75400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 553674 75200 555570 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 556154 75200 558200 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 558524 75200 560570 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 561230 75200 563276 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 563600 75200 565646 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 566230 75200 568126 75400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 579474 75200 581370 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 581954 75200 584000 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 584324 75200 586370 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 587030 75200 589076 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 589400 75200 591446 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 592030 75200 593926 75400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal5 710930 90774 711200 92670 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 93254 711200 95300 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 95624 711200 97670 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 98330 711200 100376 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 100700 711200 102746 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 103330 711200 105226 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 710930 118974 711200 120870 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 121454 711200 123500 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 123824 711200 125870 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 126530 711200 128576 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 128900 711200 130946 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 131530 711200 133426 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 710930 372774 711200 374670 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 375254 711200 377300 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 377624 711200 379670 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 380330 711200 382376 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 382700 711200 384746 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 385330 711200 387226 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 710930 400974 711200 402870 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 710930 403454 711200 405500 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 710930 405824 711200 407870 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 710930 408530 711200 410576 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 710930 410900 711200 412946 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 710930 413530 711200 415426 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal4 579474 430800 581370 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 581954 430800 584000 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 584324 430800 586370 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 587030 430800 589076 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 589400 430800 591446 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 592030 430800 593926 431000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal4 553674 430800 555570 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 556154 430800 558200 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 558524 430800 560570 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 561230 430800 563276 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 563600 430800 565646 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 566230 430800 568126 431000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal4 218274 430800 220170 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 220754 430800 222800 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 223124 430800 225170 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 225830 430800 227876 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 228200 430800 230246 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 230830 430800 232726 431000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal4 192474 430800 194370 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 194954 430800 197000 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 197324 430800 199370 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 200030 430800 202076 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 202400 430800 204446 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal4 205030 430800 206926 431000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew
flabel metal5 75200 413530 75470 415426 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 410900 75470 412946 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 408530 75470 410576 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 405824 75470 407870 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 403454 75470 405500 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 400974 75470 402870 0 FreeSans 1600 90 0 0 VDD
port 3 nsew
flabel metal5 75200 385330 75470 387226 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 382700 75470 384746 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 380330 75470 382376 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 377624 75470 379670 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 375254 75470 377300 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 372774 75470 374670 0 FreeSans 1600 90 0 0 VSS
port 4 nsew
flabel metal5 75200 131530 75470 133426 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 128900 75470 130946 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 126530 75470 128576 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 123824 75470 125870 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 121454 75470 123500 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 118974 75470 120870 0 FreeSans 1600 90 0 0 DVDD
port 1 nsew
flabel metal5 75200 103330 75470 105226 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 75200 100700 75470 102746 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 75200 98330 75470 100376 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 75200 95624 75470 97670 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 75200 93254 75470 95300 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
flabel metal5 75200 90774 75470 92670 0 FreeSans 1600 90 0 0 DVSS
port 2 nsew
<< end >>
