magic
tech gf180mcuD
magscale 1 10
timestamp 1765055688
<< metal2 >>
rect -30 15114 59 15190
rect 222 15114 232 15190
rect -30 3008 59 3084
rect 222 3008 232 3084
rect -30 2135 59 2211
rect 222 2135 232 2211
rect 0 308 59 384
rect 222 308 232 384
rect 0 120 59 196
rect 222 120 232 196
<< via2 >>
rect 59 15114 222 15190
rect 59 3008 222 3084
rect 59 2135 222 2211
rect 59 308 222 384
rect 59 120 222 196
<< metal3 >>
rect 49 15114 59 15190
rect 222 15114 303 15190
rect 49 3008 59 3084
rect 222 3008 303 3084
rect 49 2135 59 2211
rect 222 2135 303 2211
rect 192 561 252 572
rect 192 398 193 561
rect 251 398 252 561
rect 192 384 252 398
rect 49 308 59 384
rect 222 308 303 384
rect 43 120 59 196
rect 222 120 303 196
rect 73 111 131 120
rect 73 -62 131 -52
<< via3 >>
rect 193 398 251 561
rect 73 -52 131 111
<< metal4 >>
rect 72 111 132 3147
rect 72 -52 73 111
rect 131 -52 132 111
rect 192 561 252 3147
rect 192 398 193 561
rect 251 398 252 561
rect 192 75 252 398
rect 72 -62 132 -52
<< properties >>
string flatten true
<< end >>
