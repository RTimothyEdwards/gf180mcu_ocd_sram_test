magic
tech gf180mcuD
magscale 1 10
timestamp 1765074952
<< checkpaint >>
rect 528281 430815 541692 430965
<< via1 >>
rect 528281 430913 528338 430965
rect 528802 430913 528859 430965
rect 529674 430913 529731 430965
rect 529885 430913 529942 430965
rect 541343 430913 541400 430965
rect 529031 430815 529088 430867
rect 529173 430815 529230 430867
rect 541635 430815 541692 430867
<< end >>
