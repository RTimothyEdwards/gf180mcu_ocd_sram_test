magic
tech gf180mcuD
magscale 1 10
timestamp 1765133588
<< metal5 >>
rect 94032 491968 99032 496968
rect 119832 491968 124832 496968
rect 145632 491968 150632 496968
rect 171432 491968 176432 496968
rect 197232 491968 202232 496968
rect 223032 491968 228032 496968
rect 248832 491968 253832 496968
rect 274632 491968 279632 496968
rect 300432 491968 305432 496968
rect 326232 491968 331232 496968
rect 352032 491968 357032 496968
rect 377832 491968 382832 496968
rect 403632 491968 408632 496968
rect 429432 491968 434432 496968
rect 455232 491968 460232 496968
rect 481032 491968 486032 496968
rect 506832 491968 511832 496968
rect 532632 491968 537632 496968
rect 558432 491968 563432 496968
rect 584232 491968 589232 496968
rect 610032 491968 615032 496968
rect 635832 491968 640832 496968
rect 661632 491968 666632 496968
rect 687432 491968 692432 496968
rect 9200 405732 14200 410732
rect 772168 405732 777168 410732
rect 9200 377532 14200 382532
rect 772168 377532 777168 382532
rect 9200 349332 14200 354332
rect 772168 349332 777168 354332
rect 9200 321132 14200 326132
rect 772168 321132 777168 326132
rect 9200 292932 14200 297932
rect 772168 292932 777168 297932
rect 9200 264732 14200 269732
rect 772168 264732 777168 269732
rect 9200 236532 14200 241532
rect 772168 236532 777168 241532
rect 9200 208332 14200 213332
rect 772168 208332 777168 213332
rect 9200 180132 14200 185132
rect 772168 180132 777168 185132
rect 9200 151932 14200 156932
rect 772168 151932 777168 156932
rect 9200 123732 14200 128732
rect 772168 123732 777168 128732
rect 9200 95532 14200 100532
rect 772168 95532 777168 100532
rect 94032 9168 99032 14168
rect 119832 9168 124832 14168
rect 145632 9168 150632 14168
rect 171432 9168 176432 14168
rect 197232 9168 202232 14168
rect 223032 9168 228032 14168
rect 248832 9168 253832 14168
rect 274632 9168 279632 14168
rect 300432 9168 305432 14168
rect 326232 9168 331232 14168
rect 352032 9168 357032 14168
rect 377832 9168 382832 14168
rect 403632 9168 408632 14168
rect 429432 9168 434432 14168
rect 455232 9168 460232 14168
rect 481032 9168 486032 14168
rect 506832 9168 511832 14168
rect 532632 9168 537632 14168
rect 558432 9168 563432 14168
rect 584232 9168 589232 14168
rect 610032 9168 615032 14168
rect 635832 9168 640832 14168
rect 661632 9168 666632 14168
rect 687432 9168 692432 14168
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 1 5200 -1 0 274700
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_1
timestamp 1765124241
transform 0 1 5200 -1 0 302900
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_2
timestamp 1765124241
transform 0 1 5200 -1 0 359300
box -32 0 15032 70000
use gf180mcu_ocd_io__asig_5p0  gf180mcu_ocd_io__asig_5p0_3
timestamp 1765124241
transform 0 1 5200 -1 0 331100
box -32 0 15032 70000
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 1 0 682400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_1
timestamp 1765124241
transform 1 0 656600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_2
timestamp 1765124241
transform 1 0 630800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_3
timestamp 1765124241
transform 1 0 605000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_4
timestamp 1765124241
transform 1 0 450200 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_5
timestamp 1765124241
transform 1 0 398600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_6
timestamp 1765124241
transform 1 0 476000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_7
timestamp 1765124241
transform 1 0 527600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_8
timestamp 1765124241
transform 1 0 501800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_9
timestamp 1765124241
transform 1 0 424400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_10
timestamp 1765124241
transform 0 -1 781200 1 0 175100
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_11
timestamp 1765124241
transform 0 -1 781200 1 0 146900
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_12
timestamp 1765124241
transform 0 -1 781200 1 0 203300
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_13
timestamp 1765124241
transform 0 -1 781200 1 0 231500
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_14
timestamp 1765124241
transform 1 0 269600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_15
timestamp 1765124241
transform 1 0 347000 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_16
timestamp 1765124241
transform 1 0 372800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_17
timestamp 1765124241
transform 1 0 295400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_18
timestamp 1765124241
transform 1 0 321200 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_19
timestamp 1765124241
transform 1 0 243800 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_20
timestamp 1765124241
transform 1 0 140600 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_21
timestamp 1765124241
transform 1 0 166400 0 1 5200
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_22
timestamp 1765124241
transform 1 0 89000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_23
timestamp 1765124241
transform 1 0 140600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_24
timestamp 1765124241
transform 1 0 166400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_25
timestamp 1765124241
transform 1 0 114800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_26
timestamp 1765124241
transform 1 0 372800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_27
timestamp 1765124241
transform 1 0 295400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_28
timestamp 1765124241
transform 1 0 347000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_29
timestamp 1765124241
transform 1 0 243800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_30
timestamp 1765124241
transform 1 0 269600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_31
timestamp 1765124241
transform 1 0 321200 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_32
timestamp 1765124241
transform 0 -1 781200 1 0 287900
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_33
timestamp 1765124241
transform 0 -1 781200 1 0 259700
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_34
timestamp 1765124241
transform 0 -1 781200 1 0 316100
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_35
timestamp 1765124241
transform 0 -1 781200 1 0 344300
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_36
timestamp 1765124241
transform 1 0 501800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_37
timestamp 1765124241
transform 1 0 476000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_38
timestamp 1765124241
transform 1 0 424400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_39
timestamp 1765124241
transform 1 0 450200 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_40
timestamp 1765124241
transform 1 0 398600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_41
timestamp 1765124241
transform 1 0 527600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_42
timestamp 1765124241
transform 1 0 630800 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_43
timestamp 1765124241
transform 1 0 656600 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_44
timestamp 1765124241
transform 1 0 682400 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_45
timestamp 1765124241
transform 1 0 605000 0 -1 501000
box -32 0 15032 70001
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform -1 0 781200 0 1 5200
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_1
timestamp 1765124241
transform 1 0 5200 0 1 5200
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_2
timestamp 1765124241
transform 1 0 5200 0 -1 501000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  gf180mcu_ocd_io__cor_3
timestamp 1765124241
transform -1 0 781200 0 -1 501000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_1 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 1 0 579200 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_3
timestamp 1765124241
transform 0 1 5200 -1 0 133700
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_5
timestamp 1765124241
transform 1 0 218000 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  gf180mcu_ocd_io__dvdd_6
timestamp 1765124241
transform 0 -1 781200 1 0 400700
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_1 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 1 0 553400 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_2
timestamp 1765124241
transform 0 1 5200 -1 0 105500
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_5
timestamp 1765124241
transform 1 0 192200 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  gf180mcu_ocd_io__dvss_7
timestamp 1765124241
transform 0 -1 781200 1 0 372500
box -32 0 15032 70000
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 118500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_1
timestamp 1765124241
transform 0 -1 781200 1 0 90200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_2
timestamp 1765124241
transform 1 0 656200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_3
timestamp 1765124241
transform 1 0 656400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_4
timestamp 1765124241
transform 1 0 681600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_5
timestamp 1765124241
transform 1 0 681800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_6
timestamp 1765124241
transform 1 0 682000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_7
timestamp 1765124241
transform 1 0 682200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_8
timestamp 1765124241
transform 1 0 709400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_9
timestamp 1765124241
transform 1 0 709600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_10
timestamp 1765124241
transform 1 0 709800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_11
timestamp 1765124241
transform 1 0 710000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_12
timestamp 1765124241
transform 1 0 656000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_13
timestamp 1765124241
transform 1 0 604200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_14
timestamp 1765124241
transform 1 0 604400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_15
timestamp 1765124241
transform 1 0 604600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_16
timestamp 1765124241
transform 1 0 604800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_17
timestamp 1765124241
transform 1 0 630000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_18
timestamp 1765124241
transform 1 0 630200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_19
timestamp 1765124241
transform 1 0 630400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_20
timestamp 1765124241
transform 1 0 630600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_21
timestamp 1765124241
transform 1 0 655800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_22
timestamp 1765124241
transform 1 0 449600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_23
timestamp 1765124241
transform 1 0 449400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_24
timestamp 1765124241
transform 1 0 424200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_25
timestamp 1765124241
transform 1 0 449800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_26
timestamp 1765124241
transform 1 0 423800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_27
timestamp 1765124241
transform 1 0 424000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_28
timestamp 1765124241
transform 1 0 450000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_29
timestamp 1765124241
transform 1 0 475200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_30
timestamp 1765124241
transform 1 0 475400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_31
timestamp 1765124241
transform 1 0 475600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_32
timestamp 1765124241
transform 1 0 475800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_33
timestamp 1765124241
transform 1 0 501000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_34
timestamp 1765124241
transform 1 0 501200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_35
timestamp 1765124241
transform 1 0 501400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_36
timestamp 1765124241
transform 1 0 501600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_37
timestamp 1765124241
transform 1 0 526800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_38
timestamp 1765124241
transform 1 0 423600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_39
timestamp 1765124241
transform 1 0 397800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_40
timestamp 1765124241
transform 1 0 398000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_41
timestamp 1765124241
transform 1 0 398200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_42
timestamp 1765124241
transform 1 0 398400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_43
timestamp 1765124241
transform 1 0 527000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_44
timestamp 1765124241
transform 1 0 527400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_45
timestamp 1765124241
transform 1 0 527200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_46
timestamp 1765124241
transform 1 0 552600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_47
timestamp 1765124241
transform 1 0 552800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_48
timestamp 1765124241
transform 1 0 553000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_49
timestamp 1765124241
transform 1 0 553200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_50
timestamp 1765124241
transform 1 0 578400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_51
timestamp 1765124241
transform 1 0 578600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_52
timestamp 1765124241
transform 1 0 578800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_53
timestamp 1765124241
transform 1 0 579000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_54
timestamp 1765124241
transform 0 -1 781200 1 0 146700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_55
timestamp 1765124241
transform 0 -1 781200 1 0 174900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_56
timestamp 1765124241
transform 0 -1 781200 1 0 203100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_57
timestamp 1765124241
transform 0 -1 781200 1 0 231300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_58
timestamp 1765124241
transform 1 0 268800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_59
timestamp 1765124241
transform 1 0 321000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_60
timestamp 1765124241
transform 1 0 320800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_61
timestamp 1765124241
transform 1 0 320600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_62
timestamp 1765124241
transform 1 0 320400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_63
timestamp 1765124241
transform 1 0 346200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_64
timestamp 1765124241
transform 1 0 346400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_65
timestamp 1765124241
transform 1 0 346600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_66
timestamp 1765124241
transform 1 0 346800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_67
timestamp 1765124241
transform 1 0 372000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_68
timestamp 1765124241
transform 1 0 269000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_69
timestamp 1765124241
transform 1 0 295200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_70
timestamp 1765124241
transform 1 0 372400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_71
timestamp 1765124241
transform 1 0 372600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_72
timestamp 1765124241
transform 1 0 295000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_73
timestamp 1765124241
transform 1 0 294800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_74
timestamp 1765124241
transform 1 0 294600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_75
timestamp 1765124241
transform 1 0 269400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_76
timestamp 1765124241
transform 1 0 269200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_77
timestamp 1765124241
transform 1 0 372200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_78
timestamp 1765124241
transform 1 0 217800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_79
timestamp 1765124241
transform 1 0 217200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_80
timestamp 1765124241
transform 1 0 217600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_81
timestamp 1765124241
transform 1 0 217400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_82
timestamp 1765124241
transform 1 0 243600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_83
timestamp 1765124241
transform 1 0 243400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_84
timestamp 1765124241
transform 1 0 243200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_85
timestamp 1765124241
transform 1 0 243000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_86
timestamp 1765124241
transform 0 1 5200 -1 0 118700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_87
timestamp 1765124241
transform 0 1 5200 -1 0 90400
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_88
timestamp 1765124241
transform 1 0 88200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_89
timestamp 1765124241
transform 1 0 88400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_90
timestamp 1765124241
transform 1 0 88600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_91
timestamp 1765124241
transform 1 0 88800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_92
timestamp 1765124241
transform 1 0 139800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_93
timestamp 1765124241
transform 1 0 140000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_94
timestamp 1765124241
transform 1 0 140400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_95
timestamp 1765124241
transform 1 0 165600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_96
timestamp 1765124241
transform 1 0 165800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_97
timestamp 1765124241
transform 1 0 166000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_98
timestamp 1765124241
transform 1 0 166200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_99
timestamp 1765124241
transform 1 0 191400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_100
timestamp 1765124241
transform 1 0 191600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_101
timestamp 1765124241
transform 1 0 191800 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_102
timestamp 1765124241
transform 1 0 192000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_103
timestamp 1765124241
transform 1 0 140200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_104
timestamp 1765124241
transform 1 0 114000 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_105
timestamp 1765124241
transform 1 0 114400 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_106
timestamp 1765124241
transform 1 0 114600 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_107
timestamp 1765124241
transform 1 0 114200 0 1 5200
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_108
timestamp 1765124241
transform 0 1 5200 -1 0 175100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_109
timestamp 1765124241
transform 0 1 5200 -1 0 146900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_110
timestamp 1765124241
transform 0 1 5200 -1 0 231500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_111
timestamp 1765124241
transform 0 1 5200 -1 0 203300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_112
timestamp 1765124241
transform 0 1 5200 -1 0 287900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_113
timestamp 1765124241
transform 0 1 5200 -1 0 259700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_114
timestamp 1765124241
transform 0 1 5200 -1 0 344300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_115
timestamp 1765124241
transform 0 1 5200 -1 0 372500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_116
timestamp 1765124241
transform 0 1 5200 -1 0 316100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_117
timestamp 1765124241
transform 0 1 5200 -1 0 429900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_118
timestamp 1765124241
transform 0 1 5200 -1 0 400700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_119
timestamp 1765124241
transform 1 0 165600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_120
timestamp 1765124241
transform 1 0 114400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_121
timestamp 1765124241
transform 1 0 88800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_122
timestamp 1765124241
transform 1 0 88600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_123
timestamp 1765124241
transform 1 0 88400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_124
timestamp 1765124241
transform 1 0 114600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_125
timestamp 1765124241
transform 1 0 88200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_126
timestamp 1765124241
transform 1 0 139800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_127
timestamp 1765124241
transform 1 0 140000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_128
timestamp 1765124241
transform 1 0 140200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_129
timestamp 1765124241
transform 1 0 140400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_130
timestamp 1765124241
transform 1 0 191400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_131
timestamp 1765124241
transform 1 0 191600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_132
timestamp 1765124241
transform 1 0 166200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_133
timestamp 1765124241
transform 1 0 191800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_134
timestamp 1765124241
transform 1 0 166000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_135
timestamp 1765124241
transform 1 0 165800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_136
timestamp 1765124241
transform 1 0 192000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_137
timestamp 1765124241
transform 1 0 114000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_138
timestamp 1765124241
transform 1 0 114200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_139
timestamp 1765124241
transform 1 0 321000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_140
timestamp 1765124241
transform 1 0 269000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_141
timestamp 1765124241
transform 1 0 320800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_142
timestamp 1765124241
transform 1 0 269400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_143
timestamp 1765124241
transform 1 0 294600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_144
timestamp 1765124241
transform 1 0 294800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_145
timestamp 1765124241
transform 1 0 295000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_146
timestamp 1765124241
transform 1 0 295200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_147
timestamp 1765124241
transform 1 0 320400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_148
timestamp 1765124241
transform 1 0 320600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_149
timestamp 1765124241
transform 1 0 269200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_150
timestamp 1765124241
transform 1 0 346200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_151
timestamp 1765124241
transform 1 0 243400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_152
timestamp 1765124241
transform 1 0 243200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_153
timestamp 1765124241
transform 1 0 243000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_154
timestamp 1765124241
transform 1 0 268800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_155
timestamp 1765124241
transform 1 0 217200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_156
timestamp 1765124241
transform 1 0 217800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_157
timestamp 1765124241
transform 1 0 217600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_158
timestamp 1765124241
transform 1 0 217400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_159
timestamp 1765124241
transform 1 0 243600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_160
timestamp 1765124241
transform 1 0 346400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_161
timestamp 1765124241
transform 1 0 372600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_162
timestamp 1765124241
transform 1 0 372400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_163
timestamp 1765124241
transform 1 0 372200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_164
timestamp 1765124241
transform 1 0 372000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_165
timestamp 1765124241
transform 1 0 346800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_166
timestamp 1765124241
transform 1 0 346600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_167
timestamp 1765124241
transform 0 -1 781200 1 0 287700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_168
timestamp 1765124241
transform 0 -1 781200 1 0 259500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_169
timestamp 1765124241
transform 0 -1 781200 1 0 315900
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_170
timestamp 1765124241
transform 0 -1 781200 1 0 344100
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_171
timestamp 1765124241
transform 0 -1 781200 1 0 372300
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_172
timestamp 1765124241
transform 1 0 579000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_173
timestamp 1765124241
transform 1 0 450000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_174
timestamp 1765124241
transform 1 0 449800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_175
timestamp 1765124241
transform 1 0 578400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_176
timestamp 1765124241
transform 1 0 578600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_177
timestamp 1765124241
transform 1 0 527400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_178
timestamp 1765124241
transform 1 0 527200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_179
timestamp 1765124241
transform 1 0 527000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_180
timestamp 1765124241
transform 1 0 526800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_181
timestamp 1765124241
transform 1 0 552600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_182
timestamp 1765124241
transform 1 0 501600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_183
timestamp 1765124241
transform 1 0 552800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_184
timestamp 1765124241
transform 1 0 449600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_185
timestamp 1765124241
transform 1 0 501200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_186
timestamp 1765124241
transform 1 0 501000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_187
timestamp 1765124241
transform 1 0 553000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_188
timestamp 1765124241
transform 1 0 553200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_189
timestamp 1765124241
transform 1 0 578800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_190
timestamp 1765124241
transform 1 0 475800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_191
timestamp 1765124241
transform 1 0 475600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_192
timestamp 1765124241
transform 1 0 475400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_193
timestamp 1765124241
transform 1 0 475200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_194
timestamp 1765124241
transform 1 0 501400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_195
timestamp 1765124241
transform 1 0 449400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_196
timestamp 1765124241
transform 1 0 424200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_197
timestamp 1765124241
transform 1 0 424000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_198
timestamp 1765124241
transform 1 0 423800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_199
timestamp 1765124241
transform 1 0 423600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_200
timestamp 1765124241
transform 1 0 398400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_201
timestamp 1765124241
transform 1 0 398000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_202
timestamp 1765124241
transform 1 0 397800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_203
timestamp 1765124241
transform 1 0 398200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_204
timestamp 1765124241
transform 0 -1 781200 1 0 429700
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_205
timestamp 1765124241
transform 0 -1 781200 1 0 400500
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_206
timestamp 1765124241
transform 1 0 681600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_207
timestamp 1765124241
transform 1 0 682200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_208
timestamp 1765124241
transform 1 0 682000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_209
timestamp 1765124241
transform 1 0 630000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_210
timestamp 1765124241
transform 1 0 681800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_211
timestamp 1765124241
transform 1 0 656400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_212
timestamp 1765124241
transform 1 0 709800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_213
timestamp 1765124241
transform 1 0 656200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_214
timestamp 1765124241
transform 1 0 656000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_215
timestamp 1765124241
transform 1 0 655800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_216
timestamp 1765124241
transform 1 0 604800 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_217
timestamp 1765124241
transform 1 0 604200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_218
timestamp 1765124241
transform 1 0 604400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_219
timestamp 1765124241
transform 1 0 604600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_220
timestamp 1765124241
transform 1 0 710000 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_221
timestamp 1765124241
transform 1 0 630200 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_222
timestamp 1765124241
transform 1 0 630400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_223
timestamp 1765124241
transform 1 0 709400 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_224
timestamp 1765124241
transform 1 0 630600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill1  gf180mcu_ocd_io__fill1_225
timestamp 1765124241
transform 1 0 709600 0 -1 501000
box -32 13097 232 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 117500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_1
timestamp 1765124241
transform 0 -1 781200 1 0 173900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_2
timestamp 1765124241
transform 0 -1 781200 1 0 145700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_3
timestamp 1765124241
transform 0 -1 781200 1 0 202100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_4
timestamp 1765124241
transform 0 -1 781200 1 0 230300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_5
timestamp 1765124241
transform 0 1 5200 -1 0 118500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_6
timestamp 1765124241
transform 0 1 5200 -1 0 174900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_7
timestamp 1765124241
transform 0 1 5200 -1 0 146700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_8
timestamp 1765124241
transform 0 1 5200 -1 0 203100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_9
timestamp 1765124241
transform 0 1 5200 -1 0 231300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_10
timestamp 1765124241
transform 0 1 5200 -1 0 259500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_11
timestamp 1765124241
transform 0 1 5200 -1 0 287700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_12
timestamp 1765124241
transform 0 1 5200 -1 0 372300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_13
timestamp 1765124241
transform 0 1 5200 -1 0 344100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_14
timestamp 1765124241
transform 0 1 5200 -1 0 315900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_15
timestamp 1765124241
transform 0 1 5200 -1 0 400500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_16
timestamp 1765124241
transform 0 -1 781200 1 0 258500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_17
timestamp 1765124241
transform 0 -1 781200 1 0 286700
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_18
timestamp 1765124241
transform 0 -1 781200 1 0 371300
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_19
timestamp 1765124241
transform 0 -1 781200 1 0 343100
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_20
timestamp 1765124241
transform 0 -1 781200 1 0 314900
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_21
timestamp 1765124241
transform 0 -1 781200 1 0 399500
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 115500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1
timestamp 1765124241
transform 0 -1 781200 1 0 105500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_2
timestamp 1765124241
transform 0 -1 781200 1 0 82200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_3
timestamp 1765124241
transform 0 -1 781200 1 0 107500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_4
timestamp 1765124241
transform 0 -1 781200 1 0 80200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_5
timestamp 1765124241
transform 0 -1 781200 1 0 78200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_6
timestamp 1765124241
transform 0 -1 781200 1 0 86200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_7
timestamp 1765124241
transform 0 -1 781200 1 0 76200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_8
timestamp 1765124241
transform 0 -1 781200 1 0 113500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_9
timestamp 1765124241
transform 0 -1 781200 1 0 111500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_10
timestamp 1765124241
transform 0 -1 781200 1 0 88200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_11
timestamp 1765124241
transform 0 -1 781200 1 0 84200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_12
timestamp 1765124241
transform 0 -1 781200 1 0 109500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_14
timestamp 1765124241
transform 1 0 679600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_15
timestamp 1765124241
transform 1 0 677600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_16
timestamp 1765124241
transform 1 0 675600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_17
timestamp 1765124241
transform 1 0 673600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_18
timestamp 1765124241
transform 1 0 626000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_19
timestamp 1765124241
transform 1 0 624000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_20
timestamp 1765124241
transform 1 0 628000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_21
timestamp 1765124241
transform 1 0 622000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_23
timestamp 1765124241
transform 1 0 602200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_24
timestamp 1765124241
transform 1 0 600200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_26
timestamp 1765124241
transform 1 0 598200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_27
timestamp 1765124241
transform 1 0 596200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_28
timestamp 1765124241
transform 1 0 594200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_29
timestamp 1765124241
transform 1 0 647800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_30
timestamp 1765124241
transform 1 0 649800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_31
timestamp 1765124241
transform 1 0 651800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_32
timestamp 1765124241
transform 1 0 653800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_33
timestamp 1765124241
transform 1 0 703400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_34
timestamp 1765124241
transform 1 0 705400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_35
timestamp 1765124241
transform 1 0 699400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_37
timestamp 1765124241
transform 1 0 701400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_38
timestamp 1765124241
transform 1 0 707400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_39
timestamp 1765124241
transform 1 0 568400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_40
timestamp 1765124241
transform 1 0 471200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_41
timestamp 1765124241
transform 1 0 570400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_42
timestamp 1765124241
transform 1 0 497000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_44
timestamp 1765124241
transform 1 0 550600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_45
timestamp 1765124241
transform 1 0 447400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_46
timestamp 1765124241
transform 1 0 495000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_48
timestamp 1765124241
transform 1 0 467200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_49
timestamp 1765124241
transform 1 0 469200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_50
timestamp 1765124241
transform 1 0 445400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_51
timestamp 1765124241
transform 1 0 576400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_52
timestamp 1765124241
transform 1 0 493000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_53
timestamp 1765124241
transform 1 0 473200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_55
timestamp 1765124241
transform 1 0 415600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_56
timestamp 1765124241
transform 1 0 417600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_57
timestamp 1765124241
transform 1 0 419600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_60
timestamp 1765124241
transform 1 0 524800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_61
timestamp 1765124241
transform 1 0 572400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_62
timestamp 1765124241
transform 1 0 395800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_63
timestamp 1765124241
transform 1 0 393800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_64
timestamp 1765124241
transform 1 0 520800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_66
timestamp 1765124241
transform 1 0 441400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_67
timestamp 1765124241
transform 1 0 548600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_68
timestamp 1765124241
transform 1 0 499000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_69
timestamp 1765124241
transform 1 0 443400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_70
timestamp 1765124241
transform 1 0 518800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_72
timestamp 1765124241
transform 1 0 546600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_73
timestamp 1765124241
transform 1 0 522800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_74
timestamp 1765124241
transform 1 0 421600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_75
timestamp 1765124241
transform 1 0 544600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_76
timestamp 1765124241
transform 0 -1 781200 1 0 165900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_77
timestamp 1765124241
transform 0 -1 781200 1 0 163900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_79
timestamp 1765124241
transform 0 -1 781200 1 0 141700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_80
timestamp 1765124241
transform 0 -1 781200 1 0 139700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_81
timestamp 1765124241
transform 0 -1 781200 1 0 137700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_82
timestamp 1765124241
transform 0 -1 781200 1 0 135700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_83
timestamp 1765124241
transform 0 -1 781200 1 0 133700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_84
timestamp 1765124241
transform 0 -1 781200 1 0 143700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_85
timestamp 1765124241
transform 0 -1 781200 1 0 169900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_86
timestamp 1765124241
transform 0 -1 781200 1 0 171900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_87
timestamp 1765124241
transform 0 -1 781200 1 0 167900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_88
timestamp 1765124241
transform 0 -1 781200 1 0 224300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_89
timestamp 1765124241
transform 0 -1 781200 1 0 226300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_90
timestamp 1765124241
transform 0 -1 781200 1 0 222300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_91
timestamp 1765124241
transform 0 -1 781200 1 0 220300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_92
timestamp 1765124241
transform 0 -1 781200 1 0 228300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_95
timestamp 1765124241
transform 0 -1 781200 1 0 248500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_96
timestamp 1765124241
transform 0 -1 781200 1 0 200100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_97
timestamp 1765124241
transform 0 -1 781200 1 0 198100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_98
timestamp 1765124241
transform 0 -1 781200 1 0 196100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_99
timestamp 1765124241
transform 0 -1 781200 1 0 194100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_100
timestamp 1765124241
transform 0 -1 781200 1 0 192100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_101
timestamp 1765124241
transform 0 -1 781200 1 0 250500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_104
timestamp 1765124241
transform 1 0 260800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_105
timestamp 1765124241
transform 1 0 237000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_107
timestamp 1765124241
transform 1 0 314400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_108
timestamp 1765124241
transform 1 0 312400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_109
timestamp 1765124241
transform 1 0 235000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_110
timestamp 1765124241
transform 1 0 286600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_111
timestamp 1765124241
transform 1 0 288600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_112
timestamp 1765124241
transform 1 0 290600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_114
timestamp 1765124241
transform 1 0 266800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_115
timestamp 1765124241
transform 1 0 241000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_116
timestamp 1765124241
transform 1 0 292600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_117
timestamp 1765124241
transform 1 0 264800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_118
timestamp 1765124241
transform 1 0 262800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_119
timestamp 1765124241
transform 1 0 239000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_120
timestamp 1765124241
transform 1 0 233000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_122
timestamp 1765124241
transform 1 0 366000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_123
timestamp 1765124241
transform 1 0 318400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_124
timestamp 1765124241
transform 1 0 389800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_125
timestamp 1765124241
transform 1 0 364000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_127
timestamp 1765124241
transform 1 0 211200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_128
timestamp 1765124241
transform 1 0 209200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_129
timestamp 1765124241
transform 1 0 344200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_130
timestamp 1765124241
transform 1 0 207200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_131
timestamp 1765124241
transform 1 0 342200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_132
timestamp 1765124241
transform 1 0 340200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_133
timestamp 1765124241
transform 1 0 213200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_134
timestamp 1765124241
transform 1 0 338200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_135
timestamp 1765124241
transform 1 0 368000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_136
timestamp 1765124241
transform 1 0 316400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_137
timestamp 1765124241
transform 1 0 370000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_139
timestamp 1765124241
transform 1 0 215200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_140
timestamp 1765124241
transform 0 1 5200 -1 0 82200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_141
timestamp 1765124241
transform 0 1 5200 -1 0 84200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_142
timestamp 1765124241
transform 0 1 5200 -1 0 80200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_143
timestamp 1765124241
transform 0 1 5200 -1 0 88200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_144
timestamp 1765124241
transform 0 1 5200 -1 0 86200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_145
timestamp 1765124241
transform 0 1 5200 -1 0 78200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_146
timestamp 1765124241
transform 0 1 5200 -1 0 90200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_147
timestamp 1765124241
transform 0 1 5200 -1 0 107500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_148
timestamp 1765124241
transform 0 1 5200 -1 0 109500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_149
timestamp 1765124241
transform 0 1 5200 -1 0 111500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_150
timestamp 1765124241
transform 0 1 5200 -1 0 113500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_151
timestamp 1765124241
transform 0 1 5200 -1 0 115500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_152
timestamp 1765124241
transform 0 1 5200 -1 0 117500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_153
timestamp 1765124241
transform 1 0 106000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_155
timestamp 1765124241
transform 1 0 108000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_156
timestamp 1765124241
transform 1 0 112000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_157
timestamp 1765124241
transform 1 0 110000 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_158
timestamp 1765124241
transform 1 0 163600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_159
timestamp 1765124241
transform 1 0 161600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_160
timestamp 1765124241
transform 1 0 159600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_161
timestamp 1765124241
transform 1 0 157600 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_162
timestamp 1765124241
transform 1 0 131800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_164
timestamp 1765124241
transform 1 0 86200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_165
timestamp 1765124241
transform 1 0 137800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_166
timestamp 1765124241
transform 1 0 135800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_167
timestamp 1765124241
transform 1 0 133800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_168
timestamp 1765124241
transform 1 0 187400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_169
timestamp 1765124241
transform 1 0 185400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_170
timestamp 1765124241
transform 1 0 183400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_172
timestamp 1765124241
transform 1 0 189400 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_173
timestamp 1765124241
transform 1 0 78200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_174
timestamp 1765124241
transform 1 0 76200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_175
timestamp 1765124241
transform 1 0 84200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_176
timestamp 1765124241
transform 1 0 80200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_178
timestamp 1765124241
transform 1 0 82200 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_179
timestamp 1765124241
transform 0 1 5200 -1 0 167900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_180
timestamp 1765124241
transform 0 1 5200 -1 0 169900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_181
timestamp 1765124241
transform 0 1 5200 -1 0 171900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_182
timestamp 1765124241
transform 0 1 5200 -1 0 173900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_183
timestamp 1765124241
transform 0 1 5200 -1 0 135700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_184
timestamp 1765124241
transform 0 1 5200 -1 0 165900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_185
timestamp 1765124241
transform 0 1 5200 -1 0 137700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_186
timestamp 1765124241
transform 0 1 5200 -1 0 139700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_187
timestamp 1765124241
transform 0 1 5200 -1 0 141700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_188
timestamp 1765124241
transform 0 1 5200 -1 0 143700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_189
timestamp 1765124241
transform 0 1 5200 -1 0 145700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_191
timestamp 1765124241
transform 0 1 5200 -1 0 194100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_192
timestamp 1765124241
transform 0 1 5200 -1 0 196100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_193
timestamp 1765124241
transform 0 1 5200 -1 0 226300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_194
timestamp 1765124241
transform 0 1 5200 -1 0 198100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_195
timestamp 1765124241
transform 0 1 5200 -1 0 200100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_196
timestamp 1765124241
transform 0 1 5200 -1 0 202100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_198
timestamp 1765124241
transform 0 1 5200 -1 0 222300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_199
timestamp 1765124241
transform 0 1 5200 -1 0 224300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_200
timestamp 1765124241
transform 0 1 5200 -1 0 250500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_201
timestamp 1765124241
transform 0 1 5200 -1 0 252500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_202
timestamp 1765124241
transform 0 1 5200 -1 0 228300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_203
timestamp 1765124241
transform 0 1 5200 -1 0 230300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_206
timestamp 1765124241
transform 0 1 5200 -1 0 284700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_207
timestamp 1765124241
transform 0 1 5200 -1 0 282700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_208
timestamp 1765124241
transform 0 1 5200 -1 0 280700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_209
timestamp 1765124241
transform 0 1 5200 -1 0 278700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_210
timestamp 1765124241
transform 0 1 5200 -1 0 276700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_211
timestamp 1765124241
transform 0 1 5200 -1 0 258500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_212
timestamp 1765124241
transform 0 1 5200 -1 0 256500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_213
timestamp 1765124241
transform 0 1 5200 -1 0 286700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_214
timestamp 1765124241
transform 0 1 5200 -1 0 314900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_215
timestamp 1765124241
transform 0 1 5200 -1 0 312900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_216
timestamp 1765124241
transform 0 1 5200 -1 0 310900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_217
timestamp 1765124241
transform 0 1 5200 -1 0 308900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_218
timestamp 1765124241
transform 0 1 5200 -1 0 306900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_219
timestamp 1765124241
transform 0 1 5200 -1 0 304900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_220
timestamp 1765124241
transform 0 1 5200 -1 0 333100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_221
timestamp 1765124241
transform 0 1 5200 -1 0 335100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_222
timestamp 1765124241
transform 0 1 5200 -1 0 371300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_223
timestamp 1765124241
transform 0 1 5200 -1 0 369300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_224
timestamp 1765124241
transform 0 1 5200 -1 0 367300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_225
timestamp 1765124241
transform 0 1 5200 -1 0 365300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_226
timestamp 1765124241
transform 0 1 5200 -1 0 363300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_227
timestamp 1765124241
transform 0 1 5200 -1 0 343100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_228
timestamp 1765124241
transform 0 1 5200 -1 0 341100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_229
timestamp 1765124241
transform 0 1 5200 -1 0 361300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_230
timestamp 1765124241
transform 0 1 5200 -1 0 339100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_231
timestamp 1765124241
transform 0 1 5200 -1 0 337100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_232
timestamp 1765124241
transform 0 1 5200 -1 0 423700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_233
timestamp 1765124241
transform 0 1 5200 -1 0 425700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_234
timestamp 1765124241
transform 0 1 5200 -1 0 427700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_235
timestamp 1765124241
transform 0 1 5200 -1 0 419700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_236
timestamp 1765124241
transform 0 1 5200 -1 0 429700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_237
timestamp 1765124241
transform 0 1 5200 -1 0 417700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_238
timestamp 1765124241
transform 0 1 5200 -1 0 399500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_239
timestamp 1765124241
transform 0 1 5200 -1 0 395500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_240
timestamp 1765124241
transform 0 1 5200 -1 0 393500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_241
timestamp 1765124241
transform 0 1 5200 -1 0 391500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_242
timestamp 1765124241
transform 0 1 5200 -1 0 389500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_243
timestamp 1765124241
transform 0 1 5200 -1 0 397500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_244
timestamp 1765124241
transform 0 1 5200 -1 0 421700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_245
timestamp 1765124241
transform 1 0 131800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_246
timestamp 1765124241
transform 1 0 133800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_248
timestamp 1765124241
transform 1 0 135800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_249
timestamp 1765124241
transform 1 0 76200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_250
timestamp 1765124241
transform 1 0 78200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_251
timestamp 1765124241
transform 1 0 80200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_252
timestamp 1765124241
transform 1 0 82200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_253
timestamp 1765124241
transform 1 0 84200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_254
timestamp 1765124241
transform 1 0 86200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_255
timestamp 1765124241
transform 1 0 189400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_256
timestamp 1765124241
transform 1 0 185400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_257
timestamp 1765124241
transform 1 0 183400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_259
timestamp 1765124241
transform 1 0 159600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_260
timestamp 1765124241
transform 1 0 163600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_261
timestamp 1765124241
transform 1 0 161600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_262
timestamp 1765124241
transform 1 0 187400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_263
timestamp 1765124241
transform 1 0 137800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_265
timestamp 1765124241
transform 1 0 157600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_267
timestamp 1765124241
transform 1 0 106000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_268
timestamp 1765124241
transform 1 0 108000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_269
timestamp 1765124241
transform 1 0 110000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_270
timestamp 1765124241
transform 1 0 112000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_272
timestamp 1765124241
transform 1 0 389800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_273
timestamp 1765124241
transform 1 0 266800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_274
timestamp 1765124241
transform 1 0 264800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_275
timestamp 1765124241
transform 1 0 262800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_276
timestamp 1765124241
transform 1 0 318400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_277
timestamp 1765124241
transform 1 0 316400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_278
timestamp 1765124241
transform 1 0 314400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_279
timestamp 1765124241
transform 1 0 312400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_281
timestamp 1765124241
transform 1 0 338200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_282
timestamp 1765124241
transform 1 0 292600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_283
timestamp 1765124241
transform 1 0 340200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_284
timestamp 1765124241
transform 1 0 290600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_285
timestamp 1765124241
transform 1 0 342200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_286
timestamp 1765124241
transform 1 0 344200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_288
timestamp 1765124241
transform 1 0 364000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_289
timestamp 1765124241
transform 1 0 366000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_290
timestamp 1765124241
transform 1 0 288600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_291
timestamp 1765124241
transform 1 0 368000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_292
timestamp 1765124241
transform 1 0 370000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_293
timestamp 1765124241
transform 1 0 286600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_295
timestamp 1765124241
transform 1 0 213200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_296
timestamp 1765124241
transform 1 0 211200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_297
timestamp 1765124241
transform 1 0 209200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_298
timestamp 1765124241
transform 1 0 207200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_299
timestamp 1765124241
transform 1 0 260800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_301
timestamp 1765124241
transform 1 0 241000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_302
timestamp 1765124241
transform 1 0 239000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_303
timestamp 1765124241
transform 1 0 237000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_304
timestamp 1765124241
transform 1 0 235000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_305
timestamp 1765124241
transform 1 0 233000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_306
timestamp 1765124241
transform 1 0 215200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_308
timestamp 1765124241
transform 0 -1 781200 1 0 282700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_309
timestamp 1765124241
transform 0 -1 781200 1 0 284700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10_310x
timestamp 1765133588
transform 0 -1 781200 1 0 302900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_311
timestamp 1765124241
transform 0 -1 781200 1 0 304900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_312
timestamp 1765124241
transform 0 -1 781200 1 0 306900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_313
timestamp 1765124241
transform 0 -1 781200 1 0 308900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_314
timestamp 1765124241
transform 0 -1 781200 1 0 310900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_315
timestamp 1765124241
transform 0 -1 781200 1 0 312900
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_316
timestamp 1765124241
transform 0 -1 781200 1 0 254500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_317
timestamp 1765124241
transform 0 -1 781200 1 0 256500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_319
timestamp 1765124241
transform 0 -1 781200 1 0 276700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_320
timestamp 1765124241
transform 0 -1 781200 1 0 278700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_321
timestamp 1765124241
transform 0 -1 781200 1 0 280700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_322
timestamp 1765124241
transform 0 -1 781200 1 0 361300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_324
timestamp 1765124241
transform 0 -1 781200 1 0 333100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_325
timestamp 1765124241
transform 0 -1 781200 1 0 335100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_326
timestamp 1765124241
transform 0 -1 781200 1 0 337100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_327
timestamp 1765124241
transform 0 -1 781200 1 0 369300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_328
timestamp 1765124241
transform 0 -1 781200 1 0 367300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_329
timestamp 1765124241
transform 0 -1 781200 1 0 365300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_330
timestamp 1765124241
transform 0 -1 781200 1 0 363300
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_332
timestamp 1765124241
transform 0 -1 781200 1 0 341100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_333
timestamp 1765124241
transform 0 -1 781200 1 0 339100
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_334
timestamp 1765124241
transform 1 0 393800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_335
timestamp 1765124241
transform 1 0 395800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_337
timestamp 1765124241
transform 1 0 415600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_338
timestamp 1765124241
transform 1 0 417600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_339
timestamp 1765124241
transform 1 0 419600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_340
timestamp 1765124241
transform 1 0 421600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_342
timestamp 1765124241
transform 1 0 441400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_343
timestamp 1765124241
transform 1 0 443400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_344
timestamp 1765124241
transform 1 0 447400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_346
timestamp 1765124241
transform 1 0 467200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_347
timestamp 1765124241
transform 1 0 469200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_348
timestamp 1765124241
transform 1 0 471200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_349
timestamp 1765124241
transform 1 0 473200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_351
timestamp 1765124241
transform 1 0 493000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_352
timestamp 1765124241
transform 1 0 495000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_353
timestamp 1765124241
transform 1 0 497000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_354
timestamp 1765124241
transform 1 0 499000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_356
timestamp 1765124241
transform 1 0 518800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_357
timestamp 1765124241
transform 1 0 445400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_358
timestamp 1765124241
transform 1 0 520800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_359
timestamp 1765124241
transform 1 0 522800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_360
timestamp 1765124241
transform 1 0 524800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_362
timestamp 1765124241
transform 1 0 544600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_363
timestamp 1765124241
transform 1 0 546600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_364
timestamp 1765124241
transform 1 0 548600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_365
timestamp 1765124241
transform 1 0 550600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_366
timestamp 1765124241
transform 1 0 568400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_367
timestamp 1765124241
transform 1 0 570400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_368
timestamp 1765124241
transform 1 0 574400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_369
timestamp 1765124241
transform 1 0 576400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_370
timestamp 1765124241
transform 1 0 572400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_371
timestamp 1765124241
transform 0 -1 781200 1 0 389500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_372
timestamp 1765124241
transform 0 -1 781200 1 0 391500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_373
timestamp 1765124241
transform 0 -1 781200 1 0 423700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_374
timestamp 1765124241
transform 0 -1 781200 1 0 421700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_375
timestamp 1765124241
transform 0 -1 781200 1 0 387500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_376
timestamp 1765124241
transform 0 -1 781200 1 0 417700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_377
timestamp 1765124241
transform 0 -1 781200 1 0 419700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_378
timestamp 1765124241
transform 0 -1 781200 1 0 397500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_379
timestamp 1765124241
transform 0 -1 781200 1 0 415700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_380
timestamp 1765124241
transform 0 -1 781200 1 0 395500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_381
timestamp 1765124241
transform 0 -1 781200 1 0 425700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_382
timestamp 1765124241
transform 0 -1 781200 1 0 393500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_383
timestamp 1765124241
transform 0 -1 781200 1 0 427700
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_384
timestamp 1765124241
transform 1 0 707400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_385
timestamp 1765124241
transform 1 0 705400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_386
timestamp 1765124241
transform 1 0 703400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_387
timestamp 1765124241
transform 1 0 602200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_388
timestamp 1765124241
transform 1 0 701400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_390
timestamp 1765124241
transform 1 0 622000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_391
timestamp 1765124241
transform 1 0 624000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_392
timestamp 1765124241
transform 1 0 626000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_393
timestamp 1765124241
transform 1 0 628000 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_394
timestamp 1765124241
transform 1 0 699400 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_396
timestamp 1765124241
transform 1 0 647800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_397
timestamp 1765124241
transform 1 0 649800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_398
timestamp 1765124241
transform 1 0 651800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_399
timestamp 1765124241
transform 1 0 653800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_402
timestamp 1765124241
transform 1 0 673600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_403
timestamp 1765124241
transform 1 0 675600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_404
timestamp 1765124241
transform 1 0 677600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_405
timestamp 1765124241
transform 1 0 679600 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_406
timestamp 1765124241
transform 1 0 600200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_407
timestamp 1765124241
transform 1 0 594200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_408
timestamp 1765124241
transform 1 0 596200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_409
timestamp 1765124241
transform 1 0 598200 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_410
timestamp 1765124241
transform 0 1 5200 -1 0 254500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_411
timestamp 1765124241
transform 1 0 391800 0 -1 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_412
timestamp 1765124241
transform 0 -1 781200 1 0 252500
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_413
timestamp 1765124241
transform 1 0 391800 0 1 5200
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_0
timestamp 1765133588
transform 0 -1 781200 1 0 218300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_13
timestamp 1765133588
transform 1 0 671600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_22
timestamp 1765133588
transform 1 0 620000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_25
timestamp 1765133588
transform 1 0 645800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_36
timestamp 1765133588
transform 1 0 697400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_43
timestamp 1765133588
transform 1 0 574400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_47
timestamp 1765133588
transform 1 0 465200 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_54
timestamp 1765133588
transform 1 0 491000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_58
timestamp 1765133588
transform 1 0 413600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_59
timestamp 1765133588
transform 1 0 542600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_65
timestamp 1765133588
transform 1 0 439400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_71
timestamp 1765133588
transform 1 0 516800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_78
timestamp 1765133588
transform 0 -1 781200 1 0 161900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_94
timestamp 1765133588
transform 0 -1 781200 1 0 246500
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_102
timestamp 1765133588
transform 0 -1 781200 1 0 190100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_103
timestamp 1765133588
transform 1 0 310400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_106
timestamp 1765133588
transform 1 0 258800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_113
timestamp 1765133588
transform 1 0 284600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_121
timestamp 1765133588
transform 1 0 336200 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_126
timestamp 1765133588
transform 1 0 362000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_138
timestamp 1765133588
transform 1 0 387800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_154
timestamp 1765133588
transform 1 0 104000 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_163
timestamp 1765133588
transform 1 0 155600 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_171
timestamp 1765133588
transform 1 0 181400 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_177
timestamp 1765133588
transform 1 0 129800 0 1 5200
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_190
timestamp 1765133588
transform 0 1 5200 1 0 161900
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_197
timestamp 1765133588
transform 0 1 5200 1 0 218300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_204
timestamp 1765133588
transform 0 1 5200 1 0 246500
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_205
timestamp 1765133588
transform 0 1 5200 1 0 190100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_247
timestamp 1765133588
transform 1 0 129800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_258
timestamp 1765133588
transform 1 0 181400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_264
timestamp 1765133588
transform 1 0 155600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_266
timestamp 1765133588
transform 1 0 104000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_271
timestamp 1765133588
transform 1 0 387800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_280
timestamp 1765133588
transform 1 0 284600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_287
timestamp 1765133588
transform 1 0 362000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_294
timestamp 1765133588
transform 1 0 310400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_300
timestamp 1765133588
transform 1 0 258800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_307
timestamp 1765133588
transform 1 0 336200 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_318
timestamp 1765133588
transform 0 -1 781200 1 0 274700
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_323
timestamp 1765133588
transform 0 -1 781200 1 0 359300
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_331
timestamp 1765133588
transform 0 -1 781200 1 0 331100
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_336
timestamp 1765133588
transform 1 0 413600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_341
timestamp 1765133588
transform 1 0 439400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_345
timestamp 1765133588
transform 1 0 465200 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_350
timestamp 1765133588
transform 1 0 491000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_355
timestamp 1765133588
transform 1 0 516800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_361
timestamp 1765133588
transform 1 0 542600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_389
timestamp 1765133588
transform 1 0 620000 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_395
timestamp 1765133588
transform 1 0 645800 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_400
timestamp 1765133588
transform 1 0 697400 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_401
timestamp 1765133588
transform 1 0 671600 0 -1 501000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 90460
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_1
timestamp 1765124241
transform 0 -1 781200 1 0 90480
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_2
timestamp 1765124241
transform 0 -1 781200 1 0 90400
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_3
timestamp 1765124241
transform 0 -1 781200 1 0 90420
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_4
timestamp 1765124241
transform 0 -1 781200 1 0 90440
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_5
timestamp 1765124241
transform 0 1 5200 -1 0 90480
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_6
timestamp 1765124241
transform 0 1 5200 -1 0 90440
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_7
timestamp 1765124241
transform 0 1 5200 -1 0 90420
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_8
timestamp 1765124241
transform 0 1 5200 -1 0 90460
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_9
timestamp 1765124241
transform 0 1 5200 -1 0 90500
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_10
timestamp 1765124241
transform 0 1 5200 -1 0 430000
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_11
timestamp 1765124241
transform 0 1 5200 -1 0 429920
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_12
timestamp 1765124241
transform 0 1 5200 -1 0 429940
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_13
timestamp 1765124241
transform 0 1 5200 -1 0 429960
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_14
timestamp 1765124241
transform 0 1 5200 -1 0 429980
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_15
timestamp 1765124241
transform 0 -1 781200 1 0 429900
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_16
timestamp 1765124241
transform 0 -1 781200 1 0 429920
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_17
timestamp 1765124241
transform 0 -1 781200 1 0 429940
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_18
timestamp 1765124241
transform 0 -1 781200 1 0 429960
box -32 13097 52 69968
use gf180mcu_ocd_io__fillnc  gf180mcu_ocd_io__fillnc_19
timestamp 1765124241
transform 0 -1 781200 1 0 429980
box -32 13097 52 69968
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform -1 0 129800 0 1 5200
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_1
timestamp 1765124241
transform 0 1 5200 -1 0 161900
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_2
timestamp 1765124241
transform 0 1 5200 -1 0 190100
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_3
timestamp 1765124241
transform 0 1 5200 -1 0 218300
box -32 0 15032 69970
use gf180mcu_ocd_io__in_c  gf180mcu_ocd_io__in_c_4
timestamp 1765124241
transform 0 1 5200 -1 0 246500
box -32 0 15032 69970
use gf180mcu_ocd_io__in_s  gf180mcu_ocd_io__in_s_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform -1 0 104000 0 1 5200
box -32 0 15032 69970
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 118700
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_2
timestamp 1765124241
transform 1 0 218000 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_4
timestamp 1765124241
transform 0 1 5200 -1 0 415700
box -32 0 15032 70000
use gf180mcu_ocd_io__vdd  gf180mcu_ocd_io__vdd_7
timestamp 1765124241
transform 1 0 579200 0 -1 501000
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765124241
transform 0 -1 781200 1 0 90500
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_3
timestamp 1765124241
transform 1 0 192200 0 1 5200
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_4
timestamp 1765124241
transform 0 1 5200 -1 0 387500
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  gf180mcu_ocd_io__vss_6
timestamp 1765124241
transform 1 0 553400 0 -1 501000
box -32 0 15032 70000
use horz_connects  horz_connects_0
timestamp 1765054368
transform 1 0 141090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_1
timestamp 1765054368
transform 1 0 166890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_2
timestamp 1765054368
transform 1 0 244290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_3
timestamp 1765054368
transform 1 0 270090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_4
timestamp 1765054368
transform 1 0 295890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_5
timestamp 1765054368
transform 1 0 321690 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_6
timestamp 1765054368
transform 1 0 347490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_7
timestamp 1765054368
transform 1 0 373290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_8
timestamp 1765054368
transform 1 0 399090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_9
timestamp 1765054368
transform 1 0 424890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_10
timestamp 1765054368
transform 1 0 450690 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_11
timestamp 1765054368
transform 1 0 476490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_12
timestamp 1765054368
transform 1 0 502290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_13
timestamp 1765054368
transform 1 0 528090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_14
timestamp 1765054368
transform 1 0 605490 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_15
timestamp 1765054368
transform 1 0 631290 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_16
timestamp 1765054368
transform 1 0 657090 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_17
timestamp 1765054368
transform 1 0 682890 0 1 75200
box 0 -48 15527 232
use horz_connects  horz_connects_18
timestamp 1765054368
transform 1 0 682890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_19
timestamp 1765054368
transform 1 0 657090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_20
timestamp 1765054368
transform 1 0 631290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_21
timestamp 1765054368
transform 1 0 605490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_22
timestamp 1765054368
transform 1 0 528090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_23
timestamp 1765054368
transform 1 0 502290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_24
timestamp 1765054368
transform 1 0 476490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_25
timestamp 1765054368
transform 1 0 450690 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_26
timestamp 1765054368
transform 1 0 424890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_27
timestamp 1765054368
transform 1 0 399090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_28
timestamp 1765054368
transform 1 0 373290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_29
timestamp 1765054368
transform 1 0 347490 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_30
timestamp 1765054368
transform 1 0 321690 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_31
timestamp 1765054368
transform 1 0 295890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_32
timestamp 1765054368
transform 1 0 270090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_33
timestamp 1765054368
transform 1 0 244290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_34
timestamp 1765054368
transform 1 0 166890 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_35
timestamp 1765054368
transform 1 0 141090 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_36
timestamp 1765054368
transform 1 0 115290 0 -1 431000
box 0 -48 15527 232
use horz_connects  horz_connects_37
timestamp 1765054368
transform 1 0 89490 0 -1 431000
box 0 -48 15527 232
use horz_connects_resetb  horz_connects_resetb_0
timestamp 1764982896
transform 1 0 115290 0 1 75170
box 12323 0 15527 232
use horz_connects_resetb  horz_connects_resetb_1
timestamp 1764982896
transform 1 0 89490 0 1 75170
box 12323 0 15527 232
use horz_power_connect  horz_power_connect_0
timestamp 1764102312
transform 1 0 192472 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_1
timestamp 1764102312
transform 1 0 218272 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_2
timestamp 1764102312
transform 1 0 553672 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_3
timestamp 1764102312
transform 1 0 579472 0 1 75200
box 0 0 14456 200
use horz_power_connect  horz_power_connect_4
timestamp 1764102312
transform -1 0 593928 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_5
timestamp 1764102312
transform -1 0 568128 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_6
timestamp 1764102312
transform -1 0 232728 0 -1 431000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_7
timestamp 1764102312
transform -1 0 206928 0 -1 431000
box 0 0 14456 200
use vert_connects  vert_connects_0
timestamp 1765055688
transform -1 0 711200 0 -1 162842
box 0 -67 303 15285
use vert_connects  vert_connects_1
timestamp 1765055688
transform -1 0 711200 0 -1 191042
box 0 -67 303 15285
use vert_connects  vert_connects_2
timestamp 1765055688
transform -1 0 711200 0 -1 219242
box 0 -67 303 15285
use vert_connects  vert_connects_3
timestamp 1765055688
transform -1 0 711200 0 -1 247442
box 0 -67 303 15285
use vert_connects  vert_connects_4
timestamp 1765055688
transform -1 0 711200 0 -1 275642
box 0 -67 303 15285
use vert_connects  vert_connects_5
timestamp 1765055688
transform -1 0 711200 0 -1 303842
box 0 -67 303 15285
use vert_connects  vert_connects_6
timestamp 1765055688
transform -1 0 711200 0 -1 332042
box 0 -67 303 15285
use vert_connects  vert_connects_7
timestamp 1765055688
transform -1 0 711200 0 -1 360242
box 0 -67 303 15285
use vert_connects_in_c  vert_connects_in_c_0
timestamp 1765055688
transform 1 0 75200 0 -1 191042
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_1
timestamp 1765055688
transform 1 0 75200 0 -1 162842
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_2
timestamp 1765055688
transform 1 0 75200 0 -1 219242
box -30 -62 303 15190
use vert_connects_in_c  vert_connects_in_c_3
timestamp 1765055688
transform 1 0 75200 0 -1 247442
box -30 -62 303 15190
use vert_power_connect  vert_power_connect_0
timestamp 1764982451
transform 1 0 710930 0 1 90772
box 0 0 270 14456
use vert_power_connect  vert_power_connect_1
timestamp 1764982451
transform 1 0 710930 0 1 118972
box 0 0 270 14456
use vert_power_connect  vert_power_connect_2
timestamp 1764982451
transform 1 0 710930 0 1 372772
box 0 0 270 14456
use vert_power_connect  vert_power_connect_3
timestamp 1764982451
transform 1 0 710930 0 1 400972
box 0 0 270 14456
use vert_power_connect  vert_power_connect_4
timestamp 1764982451
transform -1 0 75470 0 -1 415428
box 0 0 270 14456
use vert_power_connect  vert_power_connect_5
timestamp 1764982451
transform -1 0 75470 0 -1 387228
box 0 0 270 14456
use vert_power_connect  vert_power_connect_6
timestamp 1764982451
transform -1 0 75470 0 -1 133428
box 0 0 270 14456
use vert_power_connect  vert_power_connect_7
timestamp 1764982451
transform -1 0 75470 0 -1 105228
box 0 0 270 14456
<< labels >>
rlabel metal5 s 584232 9168 589232 14168 4 VDD
port 3 nsew
rlabel metal5 s 223032 9168 228032 14168 4 VDD
port 3 nsew
rlabel metal5 s 558432 9168 563432 14168 4 VSS
port 5 nsew
rlabel metal5 s 197232 9168 202232 14168 4 VSS
port 5 nsew
rlabel metal5 s 584232 491968 589232 496968 4 VDD
port 3 nsew
rlabel metal5 s 223032 491968 228032 496968 4 VDD
port 3 nsew
rlabel metal5 s 558432 491968 563432 496968 4 VSS
port 5 nsew
rlabel metal5 s 197232 491968 202232 496968 4 VSS
port 5 nsew
rlabel metal5 s 9200 405732 14200 410732 4 VDD
port 3 nsew
rlabel metal5 s 9200 123732 14200 128732 4 VDD
port 3 nsew
rlabel metal5 s 9200 377532 14200 382532 4 VSS
port 5 nsew
rlabel metal5 s 9200 95532 14200 100532 4 VSS
port 5 nsew
rlabel metal5 s 772168 405732 777168 410732 4 VDD
port 3 nsew
rlabel metal5 s 772168 123732 777168 128732 4 VDD
port 3 nsew
rlabel metal5 s 772168 377532 777168 382532 4 VSS
port 5 nsew
rlabel metal5 s 772168 95532 777168 100532 4 VSS
port 5 nsew
rlabel metal5 9200 349332 14200 354332 0 analog_PAD[0]
port 6 nsew
rlabel metal5 9200 321132 14200 326132 0 analog_PAD[1]
port 7 nsew
rlabel metal5 9200 292932 14200 297932 0 analog_PAD[2]
port 8 nsew
rlabel metal5 9200 264732 14200 269732 0 analog_PAD[3]
port 9 nsew
rlabel metal5 9200 236532 14200 241532 0 input_PAD[0]
port 10 nsew
rlabel metal5 9200 208332 14200 213332 0 input_PAD[1]
port 11 nsew
rlabel metal5 9200 180132 14200 185132 0 input_PAD[2]
port 12 nsew
rlabel metal5 9200 151932 14200 156932 0 input_PAD[3]
port 13 nsew
rlabel metal5 94032 9168 99032 14168 0 clk_PAD
port 14 nsew
rlabel metal5 119832 9168 124832 14168 0 rst_n_PAD
port 15 nsew
rlabel metal5 145632 9168 150632 14168 0 bidir_PAD[0]
port 16 nsew
rlabel metal5 171432 9168 176432 14168 0 bidir_PAD[1]
port 17 nsew
rlabel metal5 248832 9168 253832 14168 0 bidir_PAD[2]
port 18 nsew
rlabel metal5 274632 9168 279632 14168 0 bidir_PAD[3]
port 19 nsew
rlabel metal5 300432 9168 305432 14168 0 bidir_PAD[4]
port 20 nsew
rlabel metal5 326232 9168 331232 14168 0 bidir_PAD[5]
port 21 nsew
rlabel metal5 352032 9168 357032 14168 0 bidir_PAD[6]
port 22 nsew
rlabel metal5 377832 9168 382832 14168 0 bidir_PAD[7]
port 23 nsew
rlabel metal5 403632 9168 408632 14168 0 bidir_PAD[8]
port 24 nsew
rlabel metal5 429432 9168 434432 14168 0 bidir_PAD[9]
port 25 nsew
rlabel metal5 455232 9168 460232 14168 0 bidir_PAD[10]
port 26 nsew
rlabel metal5 481032 9168 486032 14168 0 bidir_PAD[11]
port 27 nsew
rlabel metal5 506832 9168 511832 14168 0 bidir_PAD[12]
port 28 nsew
rlabel metal5 532632 9168 537632 14168 0 bidir_PAD[13]
port 29 nsew
rlabel metal5 610032 9168 615032 14168 0 bidir_PAD[14]
port 30 nsew
rlabel metal5 635832 9168 640832 14168 0 bidir_PAD[15]
port 31 nsew
rlabel metal5 661632 9168 666632 14168 0 bidir_PAD[16]
port 32 nsew
rlabel metal5 687432 9168 692432 14168 0 bidir_PAD[17]
port 33 nsew
rlabel metal5 772168 151932 777168 156932 0 bidir_PAD[18]
port 34 nsew
rlabel metal5 772168 180132 777168 185132 0 bidir_PAD[19]
port 35 nsew
rlabel metal5 772168 208332 777168 213332 0 bidir_PAD[20]
port 36 nsew
rlabel metal5 772168 236532 777168 241532 0 bidir_PAD[21]
port 37 nsew
rlabel metal5 772168 264732 777168 269732 0 bidir_PAD[22]
port 38 nsew
rlabel metal5 772168 292932 777168 297932 0 bidir_PAD[23]
port 39 nsew
rlabel metal5 772168 321132 777168 326132 0 bidir_PAD[24]
port 40 nsew
rlabel metal5 772168 349332 777168 354332 0 bidir_PAD[25]
port 41 nsew
rlabel metal5 687432 491968 692432 496968 0 bidir_PAD[26]
port 42 nsew
rlabel metal5 661632 491968 666632 496968 0 bidir_PAD[27]
port 43 nsew
rlabel metal5 635832 491968 640832 496968 0 bidir_PAD[28]
port 44 nsew
rlabel metal5 610032 491968 615032 496968 0 bidir_PAD[29]
port 45 nsew
rlabel metal5 532632 491968 537632 496968 0 bidir_PAD[30]
port 46 nsew
rlabel metal5 506832 491968 511832 496968 0 bidir_PAD[31]
port 47 nsew
rlabel metal5 481032 491968 486032 496968 0 bidir_PAD[32]
port 48 nsew
rlabel metal5 455232 491968 460232 496968 0 bidir_PAD[33]
port 49 nsew
rlabel metal5 429432 491968 434432 496968 0 bidir_PAD[34]
port 50 nsew
rlabel metal5 403632 491968 408632 496968 0 bidir_PAD[35]
port 51 nsew
rlabel metal5 377832 491968 382832 496968 0 bidir_PAD[36]
port 52 nsew
rlabel metal5 352032 491968 357032 496968 0 bidir_PAD[37]
port 53 nsew
rlabel metal5 326232 491968 331232 496968 0 bidir_PAD[38]
port 54 nsew
rlabel metal5 300432 491968 305432 496968 0 bidir_PAD[39]
port 55 nsew
rlabel metal5 274632 491968 279632 496968 0 bidir_PAD[40]
port 56 nsew
rlabel metal5 248832 491968 253832 496968 0 bidir_PAD[41]
port 57 nsew
rlabel metal5 171432 491968 176432 496968 0 bidir_PAD[42]
port 58 nsew
rlabel metal5 145632 491968 150632 496968 0 bidir_PAD[43]
port 59 nsew
rlabel metal5 119832 491968 124832 496968 0 bidir_PAD[44]
port 60 nsew
rlabel metal5 94032 491968 99032 496968 0 bidir_PAD[45]
port 61 nsew
<< end >>
