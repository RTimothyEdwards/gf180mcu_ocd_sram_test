magic
tech gf180mcuD
magscale 1 10
timestamp 1765074470
<< checkpaint >>
rect 141282 75235 154691 75385
<< via1 >>
rect 142888 75333 142943 75385
rect 141282 75235 141337 75287
rect 141803 75235 141858 75287
rect 142032 75235 142087 75287
rect 142174 75235 142229 75287
rect 142676 75235 142731 75287
rect 154344 75235 154399 75287
rect 154491 75235 154546 75287
rect 154636 75235 154691 75287
<< end >>
