magic
tech gf180mcuD
magscale 1 5
timestamp 1765407047
<< metal1 >>
tri 0 14144 136 14280 se
rect 136 14144 544 14280
tri 544 14144 680 14280 sw
tri 680 14144 816 14280 se
rect 816 14144 1224 14280
tri 1224 14144 1360 14280 sw
tri 1360 14144 1496 14280 se
rect 1496 14144 1904 14280
tri 1904 14144 2040 14280 sw
tri 2040 14144 2176 14280 se
rect 2176 14144 2584 14280
tri 2584 14144 2720 14280 sw
tri 2720 14144 2856 14280 se
rect 2856 14144 3264 14280
tri 3264 14144 3400 14280 sw
tri 3400 14144 3536 14280 se
rect 3536 14144 3944 14280
tri 3944 14144 4080 14280 sw
tri 4080 14144 4216 14280 se
rect 4216 14144 4624 14280
tri 4624 14144 4760 14280 sw
rect 0 13736 4760 14144
tri 0 13600 136 13736 ne
tri 0 13464 136 13600 se
rect 136 13464 544 13736
tri 544 13600 680 13736 nw
tri 680 13600 816 13736 ne
rect 816 13600 1224 13736
tri 1224 13600 1360 13736 nw
tri 1360 13600 1496 13736 ne
rect 1496 13600 1904 13736
tri 1904 13600 2040 13736 nw
tri 2040 13600 2176 13736 ne
rect 2176 13600 2584 13736
tri 2584 13600 2720 13736 nw
tri 2720 13600 2856 13736 ne
rect 2856 13600 3264 13736
tri 3264 13600 3400 13736 nw
tri 3400 13600 3536 13736 ne
rect 3536 13600 3944 13736
tri 3944 13600 4080 13736 nw
tri 4080 13600 4216 13736 ne
tri 544 13464 680 13600 sw
rect 0 13056 680 13464
tri 0 12920 136 13056 ne
tri 0 12784 136 12920 se
rect 136 12784 544 13056
tri 544 12920 680 13056 nw
tri 4080 13464 4216 13600 se
rect 4216 13464 4624 13736
tri 4624 13600 4760 13736 nw
tri 6120 14144 6256 14280 se
rect 6256 14144 6664 14280
tri 6664 14144 6800 14280 sw
tri 6800 14144 6936 14280 se
rect 6936 14144 7344 14280
tri 7344 14144 7480 14280 sw
rect 6120 13736 7480 14144
tri 6120 13600 6256 13736 ne
rect 6256 13600 6664 13736
tri 6664 13600 6800 13736 nw
tri 6800 13600 6936 13736 ne
tri 4624 13464 4760 13600 sw
rect 4080 13056 4760 13464
tri 4080 12920 4216 13056 ne
tri 544 12784 680 12920 sw
rect 0 12376 680 12784
tri 0 12240 136 12376 ne
tri 0 12104 136 12240 se
rect 136 12104 544 12376
tri 544 12240 680 12376 nw
tri 544 12104 680 12240 sw
rect 0 11696 680 12104
tri 0 11560 136 11696 ne
tri 0 11424 136 11560 se
rect 136 11424 544 11696
tri 544 11560 680 11696 nw
tri 544 11424 680 11560 sw
rect 0 11016 680 11424
tri 0 10880 136 11016 ne
tri 0 10744 136 10880 se
rect 136 10744 544 11016
tri 544 10880 680 11016 nw
tri 1360 12784 1496 12920 se
rect 1496 12784 1904 12920
tri 1904 12784 2040 12920 sw
tri 2040 12784 2176 12920 se
rect 2176 12784 2584 12920
tri 2584 12784 2720 12920 sw
tri 2720 12784 2856 12920 se
rect 2856 12784 3264 12920
tri 3264 12784 3400 12920 sw
rect 1360 12376 3400 12784
tri 1360 12240 1496 12376 ne
tri 1360 12104 1496 12240 se
rect 1496 12104 1904 12376
tri 1904 12240 2040 12376 nw
tri 2040 12240 2176 12376 ne
tri 1904 12104 2040 12240 sw
tri 2040 12104 2176 12240 se
rect 2176 12104 2584 12376
tri 2584 12240 2720 12376 nw
tri 2720 12240 2856 12376 ne
tri 2584 12104 2720 12240 sw
tri 2720 12104 2856 12240 se
rect 2856 12104 3264 12376
tri 3264 12240 3400 12376 nw
tri 3264 12104 3400 12240 sw
rect 1360 11696 3400 12104
tri 1360 11560 1496 11696 ne
tri 1360 11424 1496 11560 se
rect 1496 11424 1904 11696
tri 1904 11560 2040 11696 nw
tri 2040 11560 2176 11696 ne
tri 1904 11424 2040 11560 sw
tri 2040 11424 2176 11560 se
rect 2176 11424 2584 11696
tri 2584 11560 2720 11696 nw
tri 2720 11560 2856 11696 ne
tri 2584 11424 2720 11560 sw
tri 2720 11424 2856 11560 se
rect 2856 11424 3264 11696
tri 3264 11560 3400 11696 nw
tri 3264 11424 3400 11560 sw
rect 1360 11016 3400 11424
tri 1360 10880 1496 11016 ne
rect 1496 10880 1904 11016
tri 1904 10880 2040 11016 nw
tri 2040 10880 2176 11016 ne
rect 2176 10880 2584 11016
tri 2584 10880 2720 11016 nw
tri 2720 10880 2856 11016 ne
rect 2856 10880 3264 11016
tri 3264 10880 3400 11016 nw
tri 4080 12784 4216 12920 se
rect 4216 12784 4624 13056
tri 4624 12920 4760 13056 nw
tri 6800 13464 6936 13600 se
rect 6936 13464 7344 13736
tri 7344 13600 7480 13736 nw
tri 8160 14144 8296 14280 se
rect 8296 14144 8704 14280
tri 8704 14144 8840 14280 sw
rect 8160 13736 8840 14144
tri 8160 13600 8296 13736 ne
rect 8296 13600 8704 13736
tri 8704 13600 8840 13736 nw
tri 9520 14144 9656 14280 se
rect 9656 14144 10064 14280
tri 10064 14144 10200 14280 sw
tri 10200 14144 10336 14280 se
rect 10336 14144 10744 14280
tri 10744 14144 10880 14280 sw
tri 10880 14144 11016 14280 se
rect 11016 14144 11424 14280
tri 11424 14144 11560 14280 sw
tri 11560 14144 11696 14280 se
rect 11696 14144 12104 14280
tri 12104 14144 12240 14280 sw
tri 12240 14144 12376 14280 se
rect 12376 14144 12784 14280
tri 12784 14144 12920 14280 sw
tri 12920 14144 13056 14280 se
rect 13056 14144 13464 14280
tri 13464 14144 13600 14280 sw
tri 13600 14144 13736 14280 se
rect 13736 14144 14144 14280
tri 14144 14144 14280 14280 sw
rect 9520 13736 14280 14144
tri 9520 13600 9656 13736 ne
tri 7344 13464 7480 13600 sw
tri 7480 13464 7616 13600 se
rect 7616 13464 8024 13600
tri 8024 13464 8160 13600 sw
rect 6800 13056 8160 13464
tri 6800 12920 6936 13056 ne
rect 6936 12920 7344 13056
tri 7344 12920 7480 13056 nw
tri 7480 12920 7616 13056 ne
tri 4624 12784 4760 12920 sw
rect 4080 12376 4760 12784
tri 4080 12240 4216 12376 ne
tri 4080 12104 4216 12240 se
rect 4216 12104 4624 12376
tri 4624 12240 4760 12376 nw
tri 7480 12784 7616 12920 se
rect 7616 12784 8024 13056
tri 8024 12920 8160 13056 nw
tri 9520 13464 9656 13600 se
rect 9656 13464 10064 13736
tri 10064 13600 10200 13736 nw
tri 10200 13600 10336 13736 ne
rect 10336 13600 10744 13736
tri 10744 13600 10880 13736 nw
tri 10880 13600 11016 13736 ne
rect 11016 13600 11424 13736
tri 11424 13600 11560 13736 nw
tri 11560 13600 11696 13736 ne
rect 11696 13600 12104 13736
tri 12104 13600 12240 13736 nw
tri 12240 13600 12376 13736 ne
rect 12376 13600 12784 13736
tri 12784 13600 12920 13736 nw
tri 12920 13600 13056 13736 ne
rect 13056 13600 13464 13736
tri 13464 13600 13600 13736 nw
tri 13600 13600 13736 13736 ne
tri 10064 13464 10200 13600 sw
rect 9520 13056 10200 13464
tri 9520 12920 9656 13056 ne
tri 8024 12784 8160 12920 sw
tri 8160 12784 8296 12920 se
rect 8296 12784 8704 12920
tri 8704 12784 8840 12920 sw
rect 7480 12376 8840 12784
tri 7480 12240 7616 12376 ne
tri 4624 12104 4760 12240 sw
rect 4080 11696 4760 12104
tri 4080 11560 4216 11696 ne
tri 4080 11424 4216 11560 se
rect 4216 11424 4624 11696
tri 4624 11560 4760 11696 nw
tri 6120 12104 6256 12240 se
rect 6256 12104 6664 12240
tri 6664 12104 6800 12240 sw
rect 6120 11696 6800 12104
tri 6120 11560 6256 11696 ne
tri 4624 11424 4760 11560 sw
rect 4080 11016 4760 11424
tri 4080 10880 4216 11016 ne
tri 544 10744 680 10880 sw
rect 0 10336 680 10744
tri 0 10200 136 10336 ne
tri 0 10064 136 10200 se
rect 136 10064 544 10336
tri 544 10200 680 10336 nw
tri 4080 10744 4216 10880 se
rect 4216 10744 4624 11016
tri 4624 10880 4760 11016 nw
tri 5440 11424 5576 11560 se
rect 5576 11424 5984 11560
tri 5984 11424 6120 11560 sw
tri 6120 11424 6256 11560 se
rect 6256 11424 6664 11696
tri 6664 11560 6800 11696 nw
tri 7480 12104 7616 12240 se
rect 7616 12104 8024 12376
tri 8024 12240 8160 12376 nw
tri 8160 12240 8296 12376 ne
tri 8024 12104 8160 12240 sw
tri 8160 12104 8296 12240 se
rect 8296 12104 8704 12376
tri 8704 12240 8840 12376 nw
tri 8704 12104 8840 12240 sw
rect 7480 11696 8840 12104
tri 7480 11560 7616 11696 ne
rect 7616 11560 8024 11696
tri 8024 11560 8160 11696 nw
tri 8160 11560 8296 11696 ne
rect 8296 11560 8704 11696
tri 8704 11560 8840 11696 nw
tri 9520 12784 9656 12920 se
rect 9656 12784 10064 13056
tri 10064 12920 10200 13056 nw
tri 13600 13464 13736 13600 se
rect 13736 13464 14144 13736
tri 14144 13600 14280 13736 nw
tri 14144 13464 14280 13600 sw
rect 13600 13056 14280 13464
tri 13600 12920 13736 13056 ne
tri 10064 12784 10200 12920 sw
rect 9520 12376 10200 12784
tri 9520 12240 9656 12376 ne
tri 9520 12104 9656 12240 se
rect 9656 12104 10064 12376
tri 10064 12240 10200 12376 nw
tri 10064 12104 10200 12240 sw
rect 9520 11696 10200 12104
tri 9520 11560 9656 11696 ne
tri 6664 11424 6800 11560 sw
rect 5440 11016 6800 11424
tri 5440 10880 5576 11016 ne
rect 5576 10880 5984 11016
tri 5984 10880 6120 11016 nw
tri 6120 10880 6256 11016 ne
tri 4624 10744 4760 10880 sw
rect 4080 10336 4760 10744
tri 4080 10200 4216 10336 ne
tri 544 10064 680 10200 sw
tri 680 10064 816 10200 se
rect 816 10064 1224 10200
tri 1224 10064 1360 10200 sw
tri 1360 10064 1496 10200 se
rect 1496 10064 1904 10200
tri 1904 10064 2040 10200 sw
tri 2040 10064 2176 10200 se
rect 2176 10064 2584 10200
tri 2584 10064 2720 10200 sw
tri 2720 10064 2856 10200 se
rect 2856 10064 3264 10200
tri 3264 10064 3400 10200 sw
tri 3400 10064 3536 10200 se
rect 3536 10064 3944 10200
tri 3944 10064 4080 10200 sw
tri 4080 10064 4216 10200 se
rect 4216 10064 4624 10336
tri 4624 10200 4760 10336 nw
tri 6120 10744 6256 10880 se
rect 6256 10744 6664 11016
tri 6664 10880 6800 11016 nw
tri 9520 11424 9656 11560 se
rect 9656 11424 10064 11696
tri 10064 11560 10200 11696 nw
tri 10064 11424 10200 11560 sw
rect 9520 11016 10200 11424
tri 9520 10880 9656 11016 ne
tri 6664 10744 6800 10880 sw
tri 6800 10744 6936 10880 se
rect 6936 10744 7344 10880
tri 7344 10744 7480 10880 sw
rect 6120 10336 7480 10744
tri 6120 10200 6256 10336 ne
rect 6256 10200 6664 10336
tri 6664 10200 6800 10336 nw
tri 6800 10200 6936 10336 ne
tri 4624 10064 4760 10200 sw
rect 0 9656 4760 10064
tri 0 9520 136 9656 ne
rect 136 9520 544 9656
tri 544 9520 680 9656 nw
tri 680 9520 816 9656 ne
rect 816 9520 1224 9656
tri 1224 9520 1360 9656 nw
tri 1360 9520 1496 9656 ne
rect 1496 9520 1904 9656
tri 1904 9520 2040 9656 nw
tri 2040 9520 2176 9656 ne
rect 2176 9520 2584 9656
tri 2584 9520 2720 9656 nw
tri 2720 9520 2856 9656 ne
rect 2856 9520 3264 9656
tri 3264 9520 3400 9656 nw
tri 3400 9520 3536 9656 ne
rect 3536 9520 3944 9656
tri 3944 9520 4080 9656 nw
tri 4080 9520 4216 9656 ne
rect 4216 9520 4624 9656
tri 4624 9520 4760 9656 nw
tri 5440 10064 5576 10200 se
rect 5576 10064 5984 10200
tri 5984 10064 6120 10200 sw
rect 5440 9656 6120 10064
tri 5440 9520 5576 9656 ne
tri 5440 9384 5576 9520 se
rect 5576 9384 5984 9656
tri 5984 9520 6120 9656 nw
tri 6800 10064 6936 10200 se
rect 6936 10064 7344 10336
tri 7344 10200 7480 10336 nw
tri 7344 10064 7480 10200 sw
rect 6800 9656 7480 10064
tri 6800 9520 6936 9656 ne
tri 5984 9384 6120 9520 sw
tri 6120 9384 6256 9520 se
rect 6256 9384 6664 9520
tri 6664 9384 6800 9520 sw
tri 6800 9384 6936 9520 se
rect 6936 9384 7344 9656
tri 7344 9520 7480 9656 nw
tri 8160 10744 8296 10880 se
rect 8296 10744 8704 10880
tri 8704 10744 8840 10880 sw
rect 8160 10336 8840 10744
tri 8160 10200 8296 10336 ne
tri 8160 10064 8296 10200 se
rect 8296 10064 8704 10336
tri 8704 10200 8840 10336 nw
tri 8704 10064 8840 10200 sw
rect 8160 9656 8840 10064
tri 8160 9520 8296 9656 ne
rect 8296 9520 8704 9656
tri 8704 9520 8840 9656 nw
tri 9520 10744 9656 10880 se
rect 9656 10744 10064 11016
tri 10064 10880 10200 11016 nw
tri 10880 12784 11016 12920 se
rect 11016 12784 11424 12920
tri 11424 12784 11560 12920 sw
tri 11560 12784 11696 12920 se
rect 11696 12784 12104 12920
tri 12104 12784 12240 12920 sw
tri 12240 12784 12376 12920 se
rect 12376 12784 12784 12920
tri 12784 12784 12920 12920 sw
rect 10880 12376 12920 12784
tri 10880 12240 11016 12376 ne
tri 10880 12104 11016 12240 se
rect 11016 12104 11424 12376
tri 11424 12240 11560 12376 nw
tri 11560 12240 11696 12376 ne
tri 11424 12104 11560 12240 sw
tri 11560 12104 11696 12240 se
rect 11696 12104 12104 12376
tri 12104 12240 12240 12376 nw
tri 12240 12240 12376 12376 ne
tri 12104 12104 12240 12240 sw
tri 12240 12104 12376 12240 se
rect 12376 12104 12784 12376
tri 12784 12240 12920 12376 nw
tri 12784 12104 12920 12240 sw
rect 10880 11696 12920 12104
tri 10880 11560 11016 11696 ne
tri 10880 11424 11016 11560 se
rect 11016 11424 11424 11696
tri 11424 11560 11560 11696 nw
tri 11560 11560 11696 11696 ne
tri 11424 11424 11560 11560 sw
tri 11560 11424 11696 11560 se
rect 11696 11424 12104 11696
tri 12104 11560 12240 11696 nw
tri 12240 11560 12376 11696 ne
tri 12104 11424 12240 11560 sw
tri 12240 11424 12376 11560 se
rect 12376 11424 12784 11696
tri 12784 11560 12920 11696 nw
tri 12784 11424 12920 11560 sw
rect 10880 11016 12920 11424
tri 10880 10880 11016 11016 ne
rect 11016 10880 11424 11016
tri 11424 10880 11560 11016 nw
tri 11560 10880 11696 11016 ne
rect 11696 10880 12104 11016
tri 12104 10880 12240 11016 nw
tri 12240 10880 12376 11016 ne
rect 12376 10880 12784 11016
tri 12784 10880 12920 11016 nw
tri 13600 12784 13736 12920 se
rect 13736 12784 14144 13056
tri 14144 12920 14280 13056 nw
tri 14144 12784 14280 12920 sw
rect 13600 12376 14280 12784
tri 13600 12240 13736 12376 ne
tri 13600 12104 13736 12240 se
rect 13736 12104 14144 12376
tri 14144 12240 14280 12376 nw
tri 14144 12104 14280 12240 sw
rect 13600 11696 14280 12104
tri 13600 11560 13736 11696 ne
tri 13600 11424 13736 11560 se
rect 13736 11424 14144 11696
tri 14144 11560 14280 11696 nw
tri 14144 11424 14280 11560 sw
rect 13600 11016 14280 11424
tri 13600 10880 13736 11016 ne
tri 10064 10744 10200 10880 sw
rect 9520 10336 10200 10744
tri 9520 10200 9656 10336 ne
tri 9520 10064 9656 10200 se
rect 9656 10064 10064 10336
tri 10064 10200 10200 10336 nw
tri 13600 10744 13736 10880 se
rect 13736 10744 14144 11016
tri 14144 10880 14280 11016 nw
tri 14144 10744 14280 10880 sw
rect 13600 10336 14280 10744
tri 13600 10200 13736 10336 ne
tri 10064 10064 10200 10200 sw
tri 10200 10064 10336 10200 se
rect 10336 10064 10744 10200
tri 10744 10064 10880 10200 sw
tri 10880 10064 11016 10200 se
rect 11016 10064 11424 10200
tri 11424 10064 11560 10200 sw
tri 11560 10064 11696 10200 se
rect 11696 10064 12104 10200
tri 12104 10064 12240 10200 sw
tri 12240 10064 12376 10200 se
rect 12376 10064 12784 10200
tri 12784 10064 12920 10200 sw
tri 12920 10064 13056 10200 se
rect 13056 10064 13464 10200
tri 13464 10064 13600 10200 sw
tri 13600 10064 13736 10200 se
rect 13736 10064 14144 10336
tri 14144 10200 14280 10336 nw
tri 14144 10064 14280 10200 sw
rect 9520 9656 14280 10064
tri 9520 9520 9656 9656 ne
rect 9656 9520 10064 9656
tri 10064 9520 10200 9656 nw
tri 10200 9520 10336 9656 ne
rect 10336 9520 10744 9656
tri 10744 9520 10880 9656 nw
tri 10880 9520 11016 9656 ne
rect 11016 9520 11424 9656
tri 11424 9520 11560 9656 nw
tri 11560 9520 11696 9656 ne
rect 11696 9520 12104 9656
tri 12104 9520 12240 9656 nw
tri 12240 9520 12376 9656 ne
rect 12376 9520 12784 9656
tri 12784 9520 12920 9656 nw
tri 12920 9520 13056 9656 ne
rect 13056 9520 13464 9656
tri 13464 9520 13600 9656 nw
tri 13600 9520 13736 9656 ne
rect 13736 9520 14144 9656
tri 14144 9520 14280 9656 nw
tri 7344 9384 7480 9520 sw
rect 5440 8976 7480 9384
tri 5440 8840 5576 8976 ne
tri 1360 8704 1496 8840 se
rect 1496 8704 1904 8840
tri 1904 8704 2040 8840 sw
tri 2040 8704 2176 8840 se
rect 2176 8704 2584 8840
tri 2584 8704 2720 8840 sw
rect 1360 8296 2720 8704
tri 1360 8160 1496 8296 ne
tri 1360 8024 1496 8160 se
rect 1496 8024 1904 8296
tri 1904 8160 2040 8296 nw
tri 2040 8160 2176 8296 ne
tri 1904 8024 2040 8160 sw
tri 2040 8024 2176 8160 se
rect 2176 8024 2584 8296
tri 2584 8160 2720 8296 nw
tri 4080 8704 4216 8840 se
rect 4216 8704 4624 8840
tri 4624 8704 4760 8840 sw
tri 4760 8704 4896 8840 se
rect 4896 8704 5304 8840
tri 5304 8704 5440 8840 sw
tri 5440 8704 5576 8840 se
rect 5576 8704 5984 8976
tri 5984 8840 6120 8976 nw
tri 6120 8840 6256 8976 ne
tri 5984 8704 6120 8840 sw
tri 6120 8704 6256 8840 se
rect 6256 8704 6664 8976
tri 6664 8840 6800 8976 nw
tri 6800 8840 6936 8976 ne
rect 6936 8840 7344 8976
tri 7344 8840 7480 8976 nw
tri 6664 8704 6800 8840 sw
rect 4080 8296 6800 8704
tri 4080 8160 4216 8296 ne
rect 4216 8160 4624 8296
tri 4624 8160 4760 8296 nw
tri 4760 8160 4896 8296 ne
tri 2584 8024 2720 8160 sw
rect 1360 7616 2720 8024
tri 1360 7480 1496 7616 ne
tri 0 7344 136 7480 se
rect 136 7344 544 7480
tri 544 7344 680 7480 sw
tri 680 7344 816 7480 se
rect 816 7344 1224 7480
tri 1224 7344 1360 7480 sw
tri 1360 7344 1496 7480 se
rect 1496 7344 1904 7616
tri 1904 7480 2040 7616 nw
tri 2040 7480 2176 7616 ne
tri 1904 7344 2040 7480 sw
tri 2040 7344 2176 7480 se
rect 2176 7344 2584 7616
tri 2584 7480 2720 7616 nw
tri 4760 8024 4896 8160 se
rect 4896 8024 5304 8296
tri 5304 8160 5440 8296 nw
tri 5440 8160 5576 8296 ne
tri 5304 8024 5440 8160 sw
tri 5440 8024 5576 8160 se
rect 5576 8024 5984 8296
tri 5984 8160 6120 8296 nw
tri 6120 8160 6256 8296 ne
tri 5984 8024 6120 8160 sw
tri 6120 8024 6256 8160 se
rect 6256 8024 6664 8296
tri 6664 8160 6800 8296 nw
tri 7480 8704 7616 8840 se
rect 7616 8704 8024 8840
tri 8024 8704 8160 8840 sw
rect 7480 8296 8160 8704
tri 7480 8160 7616 8296 ne
rect 7616 8160 8024 8296
tri 8024 8160 8160 8296 nw
tri 8840 8704 8976 8840 se
rect 8976 8704 9384 8840
tri 9384 8704 9520 8840 sw
tri 9520 8704 9656 8840 se
rect 9656 8704 10064 8840
tri 10064 8704 10200 8840 sw
rect 8840 8296 10200 8704
tri 8840 8160 8976 8296 ne
tri 6664 8024 6800 8160 sw
tri 6800 8024 6936 8160 se
rect 6936 8024 7344 8160
tri 7344 8024 7480 8160 sw
rect 4760 7616 7480 8024
tri 4760 7480 4896 7616 ne
tri 2584 7344 2720 7480 sw
tri 2720 7344 2856 7480 se
rect 2856 7344 3264 7480
tri 3264 7344 3400 7480 sw
tri 3400 7344 3536 7480 se
rect 3536 7344 3944 7480
tri 3944 7344 4080 7480 sw
tri 4080 7344 4216 7480 se
rect 4216 7344 4624 7480
tri 4624 7344 4760 7480 sw
tri 4760 7344 4896 7480 se
rect 4896 7344 5304 7616
tri 5304 7480 5440 7616 nw
tri 5440 7480 5576 7616 ne
rect 5576 7480 5984 7616
tri 5984 7480 6120 7616 nw
tri 6120 7480 6256 7616 ne
tri 5304 7344 5440 7480 sw
rect 0 6936 5440 7344
tri 0 6800 136 6936 ne
rect 136 6800 544 6936
tri 544 6800 680 6936 nw
tri 680 6800 816 6936 ne
tri 680 6664 816 6800 se
rect 816 6664 1224 6936
tri 1224 6800 1360 6936 nw
tri 1360 6800 1496 6936 ne
tri 1224 6664 1360 6800 sw
tri 1360 6664 1496 6800 se
rect 1496 6664 1904 6936
tri 1904 6800 2040 6936 nw
tri 2040 6800 2176 6936 ne
rect 2176 6800 2584 6936
tri 2584 6800 2720 6936 nw
tri 2720 6800 2856 6936 ne
tri 1904 6664 2040 6800 sw
rect 680 6256 2040 6664
tri 680 6120 816 6256 ne
rect 816 6120 1224 6256
tri 1224 6120 1360 6256 nw
tri 1360 6120 1496 6256 ne
rect 1496 6120 1904 6256
tri 1904 6120 2040 6256 nw
tri 2720 6664 2856 6800 se
rect 2856 6664 3264 6936
tri 3264 6800 3400 6936 nw
tri 3400 6800 3536 6936 ne
rect 3536 6800 3944 6936
tri 3944 6800 4080 6936 nw
tri 4080 6800 4216 6936 ne
rect 4216 6800 4624 6936
tri 4624 6800 4760 6936 nw
tri 4760 6800 4896 6936 ne
tri 3264 6664 3400 6800 sw
rect 2720 6256 3400 6664
tri 2720 6120 2856 6256 ne
tri 0 5984 136 6120 se
rect 136 5984 544 6120
tri 544 5984 680 6120 sw
rect 0 5576 680 5984
tri 0 5440 136 5576 ne
rect 136 5440 544 5576
tri 544 5440 680 5576 nw
tri 2720 5984 2856 6120 se
rect 2856 5984 3264 6256
tri 3264 6120 3400 6256 nw
tri 4760 6664 4896 6800 se
rect 4896 6664 5304 6936
tri 5304 6800 5440 6936 nw
tri 6120 7344 6256 7480 se
rect 6256 7344 6664 7616
tri 6664 7480 6800 7616 nw
tri 6800 7480 6936 7616 ne
rect 6936 7480 7344 7616
tri 7344 7480 7480 7616 nw
tri 8840 8024 8976 8160 se
rect 8976 8024 9384 8296
tri 9384 8160 9520 8296 nw
tri 9520 8160 9656 8296 ne
rect 9656 8160 10064 8296
tri 10064 8160 10200 8296 nw
tri 10880 8704 11016 8840 se
rect 11016 8704 11424 8840
tri 11424 8704 11560 8840 sw
rect 10880 8296 11560 8704
tri 10880 8160 11016 8296 ne
rect 11016 8160 11424 8296
tri 11424 8160 11560 8296 nw
tri 9384 8024 9520 8160 sw
rect 8840 7616 9520 8024
tri 8840 7480 8976 7616 ne
tri 6664 7344 6800 7480 sw
rect 6120 6936 6800 7344
tri 6120 6800 6256 6936 ne
tri 5304 6664 5440 6800 sw
tri 5440 6664 5576 6800 se
rect 5576 6664 5984 6800
tri 5984 6664 6120 6800 sw
tri 6120 6664 6256 6800 se
rect 6256 6664 6664 6936
tri 6664 6800 6800 6936 nw
tri 6664 6664 6800 6800 sw
rect 4760 6256 6800 6664
tri 4760 6120 4896 6256 ne
rect 4896 6120 5304 6256
tri 5304 6120 5440 6256 nw
tri 5440 6120 5576 6256 ne
tri 3264 5984 3400 6120 sw
tri 3400 5984 3536 6120 se
rect 3536 5984 3944 6120
tri 3944 5984 4080 6120 sw
tri 4080 5984 4216 6120 se
rect 4216 5984 4624 6120
tri 4624 5984 4760 6120 sw
rect 2720 5576 4760 5984
tri 2720 5440 2856 5576 ne
rect 2856 5440 3264 5576
tri 3264 5440 3400 5576 nw
tri 3400 5440 3536 5576 ne
rect 3536 5440 3944 5576
tri 3944 5440 4080 5576 nw
tri 4080 5440 4216 5576 ne
rect 4216 5440 4624 5576
tri 4624 5440 4760 5576 nw
tri 5440 5984 5576 6120 se
rect 5576 5984 5984 6256
tri 5984 6120 6120 6256 nw
tri 6120 6120 6256 6256 ne
tri 5984 5984 6120 6120 sw
tri 6120 5984 6256 6120 se
rect 6256 5984 6664 6256
tri 6664 6120 6800 6256 nw
tri 6664 5984 6800 6120 sw
rect 5440 5576 6800 5984
tri 5440 5440 5576 5576 ne
tri 5440 5304 5576 5440 se
rect 5576 5304 5984 5576
tri 5984 5440 6120 5576 nw
tri 6120 5440 6256 5576 ne
rect 6256 5440 6664 5576
tri 6664 5440 6800 5576 nw
tri 7480 7344 7616 7480 se
rect 7616 7344 8024 7480
tri 8024 7344 8160 7480 sw
rect 7480 6936 8160 7344
tri 7480 6800 7616 6936 ne
tri 7480 6664 7616 6800 se
rect 7616 6664 8024 6936
tri 8024 6800 8160 6936 nw
tri 8840 7344 8976 7480 se
rect 8976 7344 9384 7616
tri 9384 7480 9520 7616 nw
tri 9384 7344 9520 7480 sw
rect 8840 6936 9520 7344
tri 8840 6800 8976 6936 ne
tri 8024 6664 8160 6800 sw
tri 8160 6664 8296 6800 se
rect 8296 6664 8704 6800
tri 8704 6664 8840 6800 sw
tri 8840 6664 8976 6800 se
rect 8976 6664 9384 6936
tri 9384 6800 9520 6936 nw
tri 10200 8024 10336 8160 se
rect 10336 8024 10744 8160
tri 10744 8024 10880 8160 sw
rect 10200 7616 10880 8024
tri 10200 7480 10336 7616 ne
tri 10200 7344 10336 7480 se
rect 10336 7344 10744 7616
tri 10744 7480 10880 7616 nw
tri 12240 8024 12376 8160 se
rect 12376 8024 12784 8160
tri 12784 8024 12920 8160 sw
rect 12240 7616 12920 8024
tri 12240 7480 12376 7616 ne
rect 12376 7480 12784 7616
tri 12784 7480 12920 7616 nw
tri 10744 7344 10880 7480 sw
tri 10880 7344 11016 7480 se
rect 11016 7344 11424 7480
tri 11424 7344 11560 7480 sw
tri 11560 7344 11696 7480 se
rect 11696 7344 12104 7480
tri 12104 7344 12240 7480 sw
rect 10200 6936 12240 7344
tri 10200 6800 10336 6936 ne
rect 10336 6800 10744 6936
tri 10744 6800 10880 6936 nw
tri 10880 6800 11016 6936 ne
rect 11016 6800 11424 6936
tri 11424 6800 11560 6936 nw
tri 11560 6800 11696 6936 ne
rect 11696 6800 12104 6936
tri 12104 6800 12240 6936 nw
tri 13600 7344 13736 7480 se
rect 13736 7344 14144 7480
tri 14144 7344 14280 7480 sw
rect 13600 6936 14280 7344
tri 13600 6800 13736 6936 ne
rect 13736 6800 14144 6936
tri 14144 6800 14280 6936 nw
tri 9384 6664 9520 6800 sw
tri 9520 6664 9656 6800 se
rect 9656 6664 10064 6800
tri 10064 6664 10200 6800 sw
rect 7480 6256 10200 6664
tri 7480 6120 7616 6256 ne
tri 7480 5984 7616 6120 se
rect 7616 5984 8024 6256
tri 8024 6120 8160 6256 nw
tri 8160 6120 8296 6256 ne
tri 8024 5984 8160 6120 sw
tri 8160 5984 8296 6120 se
rect 8296 5984 8704 6256
tri 8704 6120 8840 6256 nw
tri 8840 6120 8976 6256 ne
rect 8976 6120 9384 6256
tri 9384 6120 9520 6256 nw
tri 9520 6120 9656 6256 ne
rect 9656 6120 10064 6256
tri 10064 6120 10200 6256 nw
tri 12920 6664 13056 6800 se
rect 13056 6664 13464 6800
tri 13464 6664 13600 6800 sw
rect 12920 6256 13600 6664
tri 12920 6120 13056 6256 ne
rect 13056 6120 13464 6256
tri 13464 6120 13600 6256 nw
tri 8704 5984 8840 6120 sw
rect 7480 5576 8840 5984
tri 7480 5440 7616 5576 ne
tri 5984 5304 6120 5440 sw
rect 5440 4896 6120 5304
tri 5440 4760 5576 4896 ne
tri 0 4624 136 4760 se
rect 136 4624 544 4760
tri 544 4624 680 4760 sw
tri 680 4624 816 4760 se
rect 816 4624 1224 4760
tri 1224 4624 1360 4760 sw
tri 1360 4624 1496 4760 se
rect 1496 4624 1904 4760
tri 1904 4624 2040 4760 sw
tri 2040 4624 2176 4760 se
rect 2176 4624 2584 4760
tri 2584 4624 2720 4760 sw
tri 2720 4624 2856 4760 se
rect 2856 4624 3264 4760
tri 3264 4624 3400 4760 sw
tri 3400 4624 3536 4760 se
rect 3536 4624 3944 4760
tri 3944 4624 4080 4760 sw
tri 4080 4624 4216 4760 se
rect 4216 4624 4624 4760
tri 4624 4624 4760 4760 sw
rect 0 4216 4760 4624
tri 0 4080 136 4216 ne
tri 0 3944 136 4080 se
rect 136 3944 544 4216
tri 544 4080 680 4216 nw
tri 680 4080 816 4216 ne
rect 816 4080 1224 4216
tri 1224 4080 1360 4216 nw
tri 1360 4080 1496 4216 ne
rect 1496 4080 1904 4216
tri 1904 4080 2040 4216 nw
tri 2040 4080 2176 4216 ne
rect 2176 4080 2584 4216
tri 2584 4080 2720 4216 nw
tri 2720 4080 2856 4216 ne
rect 2856 4080 3264 4216
tri 3264 4080 3400 4216 nw
tri 3400 4080 3536 4216 ne
rect 3536 4080 3944 4216
tri 3944 4080 4080 4216 nw
tri 4080 4080 4216 4216 ne
tri 544 3944 680 4080 sw
rect 0 3536 680 3944
tri 0 3400 136 3536 ne
tri 0 3264 136 3400 se
rect 136 3264 544 3536
tri 544 3400 680 3536 nw
tri 4080 3944 4216 4080 se
rect 4216 3944 4624 4216
tri 4624 4080 4760 4216 nw
tri 5440 4624 5576 4760 se
rect 5576 4624 5984 4896
tri 5984 4760 6120 4896 nw
tri 6800 5304 6936 5440 se
rect 6936 5304 7344 5440
tri 7344 5304 7480 5440 sw
tri 7480 5304 7616 5440 se
rect 7616 5304 8024 5576
tri 8024 5440 8160 5576 nw
tri 8160 5440 8296 5576 ne
tri 8024 5304 8160 5440 sw
tri 8160 5304 8296 5440 se
rect 8296 5304 8704 5576
tri 8704 5440 8840 5576 nw
tri 10880 5984 11016 6120 se
rect 11016 5984 11424 6120
tri 11424 5984 11560 6120 sw
rect 10880 5576 11560 5984
tri 10880 5440 11016 5576 ne
rect 11016 5440 11424 5576
tri 11424 5440 11560 5576 nw
tri 12240 5984 12376 6120 se
rect 12376 5984 12784 6120
tri 12784 5984 12920 6120 sw
rect 12240 5576 12920 5984
tri 12240 5440 12376 5576 ne
rect 12376 5440 12784 5576
tri 12784 5440 12920 5576 nw
tri 8704 5304 8840 5440 sw
tri 8840 5304 8976 5440 se
rect 8976 5304 9384 5440
tri 9384 5304 9520 5440 sw
rect 6800 4896 9520 5304
tri 6800 4760 6936 4896 ne
tri 5984 4624 6120 4760 sw
tri 6120 4624 6256 4760 se
rect 6256 4624 6664 4760
tri 6664 4624 6800 4760 sw
tri 6800 4624 6936 4760 se
rect 6936 4624 7344 4896
tri 7344 4760 7480 4896 nw
tri 7480 4760 7616 4896 ne
tri 7344 4624 7480 4760 sw
tri 7480 4624 7616 4760 se
rect 7616 4624 8024 4896
tri 8024 4760 8160 4896 nw
tri 8160 4760 8296 4896 ne
tri 8024 4624 8160 4760 sw
tri 8160 4624 8296 4760 se
rect 8296 4624 8704 4896
tri 8704 4760 8840 4896 nw
tri 8840 4760 8976 4896 ne
rect 8976 4760 9384 4896
tri 9384 4760 9520 4896 nw
tri 10200 5304 10336 5440 se
rect 10336 5304 10744 5440
tri 10744 5304 10880 5440 sw
rect 10200 4896 10880 5304
tri 10200 4760 10336 4896 ne
rect 10336 4760 10744 4896
tri 10744 4760 10880 4896 nw
tri 11560 5304 11696 5440 se
rect 11696 5304 12104 5440
tri 12104 5304 12240 5440 sw
rect 11560 4896 12240 5304
tri 11560 4760 11696 4896 ne
rect 11696 4760 12104 4896
tri 12104 4760 12240 4896 nw
tri 13600 5304 13736 5440 se
rect 13736 5304 14144 5440
tri 14144 5304 14280 5440 sw
rect 13600 4896 14280 5304
tri 13600 4760 13736 4896 ne
rect 13736 4760 14144 4896
tri 14144 4760 14280 4896 nw
tri 8704 4624 8840 4760 sw
rect 5440 4216 8840 4624
tri 5440 4080 5576 4216 ne
rect 5576 4080 5984 4216
tri 5984 4080 6120 4216 nw
tri 6120 4080 6256 4216 ne
rect 6256 4080 6664 4216
tri 6664 4080 6800 4216 nw
tri 6800 4080 6936 4216 ne
rect 6936 4080 7344 4216
tri 7344 4080 7480 4216 nw
tri 7480 4080 7616 4216 ne
rect 7616 4080 8024 4216
tri 8024 4080 8160 4216 nw
tri 8160 4080 8296 4216 ne
rect 8296 4080 8704 4216
tri 8704 4080 8840 4216 nw
tri 10880 4624 11016 4760 se
rect 11016 4624 11424 4760
tri 11424 4624 11560 4760 sw
rect 10880 4216 11560 4624
tri 10880 4080 11016 4216 ne
rect 11016 4080 11424 4216
tri 11424 4080 11560 4216 nw
tri 12920 4624 13056 4760 se
rect 13056 4624 13464 4760
tri 13464 4624 13600 4760 sw
rect 12920 4216 13600 4624
tri 12920 4080 13056 4216 ne
rect 13056 4080 13464 4216
tri 13464 4080 13600 4216 nw
tri 4624 3944 4760 4080 sw
rect 4080 3536 4760 3944
tri 4080 3400 4216 3536 ne
tri 544 3264 680 3400 sw
rect 0 2856 680 3264
tri 0 2720 136 2856 ne
tri 0 2584 136 2720 se
rect 136 2584 544 2856
tri 544 2720 680 2856 nw
tri 544 2584 680 2720 sw
rect 0 2176 680 2584
tri 0 2040 136 2176 ne
tri 0 1904 136 2040 se
rect 136 1904 544 2176
tri 544 2040 680 2176 nw
tri 544 1904 680 2040 sw
rect 0 1496 680 1904
tri 0 1360 136 1496 ne
tri 0 1224 136 1360 se
rect 136 1224 544 1496
tri 544 1360 680 1496 nw
tri 1360 3264 1496 3400 se
rect 1496 3264 1904 3400
tri 1904 3264 2040 3400 sw
tri 2040 3264 2176 3400 se
rect 2176 3264 2584 3400
tri 2584 3264 2720 3400 sw
tri 2720 3264 2856 3400 se
rect 2856 3264 3264 3400
tri 3264 3264 3400 3400 sw
rect 1360 2856 3400 3264
tri 1360 2720 1496 2856 ne
tri 1360 2584 1496 2720 se
rect 1496 2584 1904 2856
tri 1904 2720 2040 2856 nw
tri 2040 2720 2176 2856 ne
tri 1904 2584 2040 2720 sw
tri 2040 2584 2176 2720 se
rect 2176 2584 2584 2856
tri 2584 2720 2720 2856 nw
tri 2720 2720 2856 2856 ne
tri 2584 2584 2720 2720 sw
tri 2720 2584 2856 2720 se
rect 2856 2584 3264 2856
tri 3264 2720 3400 2856 nw
tri 3264 2584 3400 2720 sw
rect 1360 2176 3400 2584
tri 1360 2040 1496 2176 ne
tri 1360 1904 1496 2040 se
rect 1496 1904 1904 2176
tri 1904 2040 2040 2176 nw
tri 2040 2040 2176 2176 ne
tri 1904 1904 2040 2040 sw
tri 2040 1904 2176 2040 se
rect 2176 1904 2584 2176
tri 2584 2040 2720 2176 nw
tri 2720 2040 2856 2176 ne
tri 2584 1904 2720 2040 sw
tri 2720 1904 2856 2040 se
rect 2856 1904 3264 2176
tri 3264 2040 3400 2176 nw
tri 3264 1904 3400 2040 sw
rect 1360 1496 3400 1904
tri 1360 1360 1496 1496 ne
rect 1496 1360 1904 1496
tri 1904 1360 2040 1496 nw
tri 2040 1360 2176 1496 ne
rect 2176 1360 2584 1496
tri 2584 1360 2720 1496 nw
tri 2720 1360 2856 1496 ne
rect 2856 1360 3264 1496
tri 3264 1360 3400 1496 nw
tri 4080 3264 4216 3400 se
rect 4216 3264 4624 3536
tri 4624 3400 4760 3536 nw
tri 9520 3944 9656 4080 se
rect 9656 3944 10064 4080
tri 10064 3944 10200 4080 sw
rect 9520 3536 10200 3944
tri 9520 3400 9656 3536 ne
tri 4624 3264 4760 3400 sw
rect 4080 2856 4760 3264
tri 4080 2720 4216 2856 ne
tri 4080 2584 4216 2720 se
rect 4216 2584 4624 2856
tri 4624 2720 4760 2856 nw
tri 6120 3264 6256 3400 se
rect 6256 3264 6664 3400
tri 6664 3264 6800 3400 sw
tri 6800 3264 6936 3400 se
rect 6936 3264 7344 3400
tri 7344 3264 7480 3400 sw
tri 7480 3264 7616 3400 se
rect 7616 3264 8024 3400
tri 8024 3264 8160 3400 sw
rect 6120 2856 8160 3264
tri 6120 2720 6256 2856 ne
rect 6256 2720 6664 2856
tri 6664 2720 6800 2856 nw
tri 6800 2720 6936 2856 ne
tri 4624 2584 4760 2720 sw
rect 4080 2176 4760 2584
tri 4080 2040 4216 2176 ne
tri 4080 1904 4216 2040 se
rect 4216 1904 4624 2176
tri 4624 2040 4760 2176 nw
tri 4624 1904 4760 2040 sw
rect 4080 1496 4760 1904
tri 4080 1360 4216 1496 ne
tri 544 1224 680 1360 sw
rect 0 816 680 1224
tri 0 680 136 816 ne
tri 0 544 136 680 se
rect 136 544 544 816
tri 544 680 680 816 nw
tri 4080 1224 4216 1360 se
rect 4216 1224 4624 1496
tri 4624 1360 4760 1496 nw
tri 5440 2584 5576 2720 se
rect 5576 2584 5984 2720
tri 5984 2584 6120 2720 sw
rect 5440 2176 6120 2584
tri 5440 2040 5576 2176 ne
tri 5440 1904 5576 2040 se
rect 5576 1904 5984 2176
tri 5984 2040 6120 2176 nw
tri 6800 2584 6936 2720 se
rect 6936 2584 7344 2856
tri 7344 2720 7480 2856 nw
tri 7480 2720 7616 2856 ne
rect 7616 2720 8024 2856
tri 8024 2720 8160 2856 nw
tri 9520 3264 9656 3400 se
rect 9656 3264 10064 3536
tri 10064 3400 10200 3536 nw
tri 12240 3944 12376 4080 se
rect 12376 3944 12784 4080
tri 12784 3944 12920 4080 sw
rect 12240 3536 12920 3944
tri 12240 3400 12376 3536 ne
rect 12376 3400 12784 3536
tri 12784 3400 12920 3536 nw
tri 13600 3944 13736 4080 se
rect 13736 3944 14144 4080
tri 14144 3944 14280 4080 sw
rect 13600 3536 14280 3944
tri 13600 3400 13736 3536 ne
tri 10064 3264 10200 3400 sw
rect 9520 2856 10200 3264
tri 9520 2720 9656 2856 ne
tri 7344 2584 7480 2720 sw
rect 6800 2176 7480 2584
tri 6800 2040 6936 2176 ne
rect 6936 2040 7344 2176
tri 7344 2040 7480 2176 nw
tri 8160 2584 8296 2720 se
rect 8296 2584 8704 2720
tri 8704 2584 8840 2720 sw
rect 8160 2176 8840 2584
tri 8160 2040 8296 2176 ne
rect 8296 2040 8704 2176
tri 8704 2040 8840 2176 nw
tri 9520 2584 9656 2720 se
rect 9656 2584 10064 2856
tri 10064 2720 10200 2856 nw
tri 11560 3264 11696 3400 se
rect 11696 3264 12104 3400
tri 12104 3264 12240 3400 sw
rect 11560 2856 12240 3264
tri 11560 2720 11696 2856 ne
rect 11696 2720 12104 2856
tri 12104 2720 12240 2856 nw
tri 13600 3264 13736 3400 se
rect 13736 3264 14144 3536
tri 14144 3400 14280 3536 nw
tri 14144 3264 14280 3400 sw
rect 13600 2856 14280 3264
tri 13600 2720 13736 2856 ne
rect 13736 2720 14144 2856
tri 14144 2720 14280 2856 nw
tri 10064 2584 10200 2720 sw
rect 9520 2176 10200 2584
tri 9520 2040 9656 2176 ne
rect 9656 2040 10064 2176
tri 10064 2040 10200 2176 nw
tri 10880 2584 11016 2720 se
rect 11016 2584 11424 2720
tri 11424 2584 11560 2720 sw
rect 10880 2176 11560 2584
tri 10880 2040 11016 2176 ne
tri 5984 1904 6120 2040 sw
rect 5440 1496 6120 1904
tri 5440 1360 5576 1496 ne
rect 5576 1360 5984 1496
tri 5984 1360 6120 1496 nw
tri 7480 1904 7616 2040 se
rect 7616 1904 8024 2040
tri 8024 1904 8160 2040 sw
rect 7480 1496 8160 1904
tri 7480 1360 7616 1496 ne
tri 4624 1224 4760 1360 sw
rect 4080 816 4760 1224
tri 4080 680 4216 816 ne
tri 544 544 680 680 sw
tri 680 544 816 680 se
rect 816 544 1224 680
tri 1224 544 1360 680 sw
tri 1360 544 1496 680 se
rect 1496 544 1904 680
tri 1904 544 2040 680 sw
tri 2040 544 2176 680 se
rect 2176 544 2584 680
tri 2584 544 2720 680 sw
tri 2720 544 2856 680 se
rect 2856 544 3264 680
tri 3264 544 3400 680 sw
tri 3400 544 3536 680 se
rect 3536 544 3944 680
tri 3944 544 4080 680 sw
tri 4080 544 4216 680 se
rect 4216 544 4624 816
tri 4624 680 4760 816 nw
tri 6120 1224 6256 1360 se
rect 6256 1224 6664 1360
tri 6664 1224 6800 1360 sw
tri 6800 1224 6936 1360 se
rect 6936 1224 7344 1360
tri 7344 1224 7480 1360 sw
tri 7480 1224 7616 1360 se
rect 7616 1224 8024 1496
tri 8024 1360 8160 1496 nw
tri 10880 1904 11016 2040 se
rect 11016 1904 11424 2176
tri 11424 2040 11560 2176 nw
tri 12920 2584 13056 2720 se
rect 13056 2584 13464 2720
tri 13464 2584 13600 2720 sw
rect 12920 2176 13600 2584
tri 12920 2040 13056 2176 ne
rect 13056 2040 13464 2176
tri 13464 2040 13600 2176 nw
tri 11424 1904 11560 2040 sw
rect 10880 1496 11560 1904
tri 10880 1360 11016 1496 ne
tri 8024 1224 8160 1360 sw
rect 6120 816 8160 1224
tri 6120 680 6256 816 ne
rect 6256 680 6664 816
tri 6664 680 6800 816 nw
tri 6800 680 6936 816 ne
rect 6936 680 7344 816
tri 7344 680 7480 816 nw
tri 7480 680 7616 816 ne
rect 7616 680 8024 816
tri 8024 680 8160 816 nw
tri 8840 1224 8976 1360 se
rect 8976 1224 9384 1360
tri 9384 1224 9520 1360 sw
rect 8840 816 9520 1224
tri 8840 680 8976 816 ne
rect 8976 680 9384 816
tri 9384 680 9520 816 nw
tri 10880 1224 11016 1360 se
rect 11016 1224 11424 1496
tri 11424 1360 11560 1496 nw
tri 12240 1904 12376 2040 se
rect 12376 1904 12784 2040
tri 12784 1904 12920 2040 sw
rect 12240 1496 12920 1904
tri 12240 1360 12376 1496 ne
rect 12376 1360 12784 1496
tri 12784 1360 12920 1496 nw
tri 11424 1224 11560 1360 sw
tri 11560 1224 11696 1360 se
rect 11696 1224 12104 1360
tri 12104 1224 12240 1360 sw
rect 10880 816 12240 1224
tri 10880 680 11016 816 ne
rect 11016 680 11424 816
tri 11424 680 11560 816 nw
tri 11560 680 11696 816 ne
rect 11696 680 12104 816
tri 12104 680 12240 816 nw
tri 12920 1224 13056 1360 se
rect 13056 1224 13464 1360
tri 13464 1224 13600 1360 sw
tri 13600 1224 13736 1360 se
rect 13736 1224 14144 1360
tri 14144 1224 14280 1360 sw
rect 12920 816 14280 1224
tri 12920 680 13056 816 ne
tri 4624 544 4760 680 sw
rect 0 136 4760 544
tri 0 0 136 136 ne
rect 136 0 544 136
tri 544 0 680 136 nw
tri 680 0 816 136 ne
rect 816 0 1224 136
tri 1224 0 1360 136 nw
tri 1360 0 1496 136 ne
rect 1496 0 1904 136
tri 1904 0 2040 136 nw
tri 2040 0 2176 136 ne
rect 2176 0 2584 136
tri 2584 0 2720 136 nw
tri 2720 0 2856 136 ne
rect 2856 0 3264 136
tri 3264 0 3400 136 nw
tri 3400 0 3536 136 ne
rect 3536 0 3944 136
tri 3944 0 4080 136 nw
tri 4080 0 4216 136 ne
rect 4216 0 4624 136
tri 4624 0 4760 136 nw
tri 8160 544 8296 680 se
rect 8296 544 8704 680
tri 8704 544 8840 680 sw
rect 8160 136 8840 544
tri 8160 0 8296 136 ne
rect 8296 0 8704 136
tri 8704 0 8840 136 nw
tri 10200 544 10336 680 se
rect 10336 544 10744 680
tri 10744 544 10880 680 sw
rect 10200 136 10880 544
tri 10200 0 10336 136 ne
rect 10336 0 10744 136
tri 10744 0 10880 136 nw
tri 12920 544 13056 680 se
rect 13056 544 13464 816
tri 13464 680 13600 816 nw
tri 13600 680 13736 816 ne
rect 13736 680 14144 816
tri 14144 680 14280 816 nw
tri 13464 544 13600 680 sw
rect 12920 136 13600 544
tri 12920 0 13056 136 ne
rect 13056 0 13464 136
tri 13464 0 13600 136 nw
<< metal2 >>
tri 0 14144 136 14280 se
rect 136 14144 544 14280
tri 544 14144 680 14280 sw
tri 680 14144 816 14280 se
rect 816 14144 1224 14280
tri 1224 14144 1360 14280 sw
tri 1360 14144 1496 14280 se
rect 1496 14144 1904 14280
tri 1904 14144 2040 14280 sw
tri 2040 14144 2176 14280 se
rect 2176 14144 2584 14280
tri 2584 14144 2720 14280 sw
tri 2720 14144 2856 14280 se
rect 2856 14144 3264 14280
tri 3264 14144 3400 14280 sw
tri 3400 14144 3536 14280 se
rect 3536 14144 3944 14280
tri 3944 14144 4080 14280 sw
tri 4080 14144 4216 14280 se
rect 4216 14144 4624 14280
tri 4624 14144 4760 14280 sw
rect 0 13736 4760 14144
tri 0 13600 136 13736 ne
tri 0 13464 136 13600 se
rect 136 13464 544 13736
tri 544 13600 680 13736 nw
tri 680 13600 816 13736 ne
rect 816 13600 1224 13736
tri 1224 13600 1360 13736 nw
tri 1360 13600 1496 13736 ne
rect 1496 13600 1904 13736
tri 1904 13600 2040 13736 nw
tri 2040 13600 2176 13736 ne
rect 2176 13600 2584 13736
tri 2584 13600 2720 13736 nw
tri 2720 13600 2856 13736 ne
rect 2856 13600 3264 13736
tri 3264 13600 3400 13736 nw
tri 3400 13600 3536 13736 ne
rect 3536 13600 3944 13736
tri 3944 13600 4080 13736 nw
tri 4080 13600 4216 13736 ne
tri 544 13464 680 13600 sw
rect 0 13056 680 13464
tri 0 12920 136 13056 ne
tri 0 12784 136 12920 se
rect 136 12784 544 13056
tri 544 12920 680 13056 nw
tri 4080 13464 4216 13600 se
rect 4216 13464 4624 13736
tri 4624 13600 4760 13736 nw
tri 6120 14144 6256 14280 se
rect 6256 14144 6664 14280
tri 6664 14144 6800 14280 sw
tri 6800 14144 6936 14280 se
rect 6936 14144 7344 14280
tri 7344 14144 7480 14280 sw
rect 6120 13736 7480 14144
tri 6120 13600 6256 13736 ne
rect 6256 13600 6664 13736
tri 6664 13600 6800 13736 nw
tri 6800 13600 6936 13736 ne
tri 4624 13464 4760 13600 sw
rect 4080 13056 4760 13464
tri 4080 12920 4216 13056 ne
tri 544 12784 680 12920 sw
rect 0 12376 680 12784
tri 0 12240 136 12376 ne
tri 0 12104 136 12240 se
rect 136 12104 544 12376
tri 544 12240 680 12376 nw
tri 544 12104 680 12240 sw
rect 0 11696 680 12104
tri 0 11560 136 11696 ne
tri 0 11424 136 11560 se
rect 136 11424 544 11696
tri 544 11560 680 11696 nw
tri 544 11424 680 11560 sw
rect 0 11016 680 11424
tri 0 10880 136 11016 ne
tri 0 10744 136 10880 se
rect 136 10744 544 11016
tri 544 10880 680 11016 nw
tri 1360 12784 1496 12920 se
rect 1496 12784 1904 12920
tri 1904 12784 2040 12920 sw
tri 2040 12784 2176 12920 se
rect 2176 12784 2584 12920
tri 2584 12784 2720 12920 sw
tri 2720 12784 2856 12920 se
rect 2856 12784 3264 12920
tri 3264 12784 3400 12920 sw
rect 1360 12376 3400 12784
tri 1360 12240 1496 12376 ne
tri 1360 12104 1496 12240 se
rect 1496 12104 1904 12376
tri 1904 12240 2040 12376 nw
tri 2040 12240 2176 12376 ne
tri 1904 12104 2040 12240 sw
tri 2040 12104 2176 12240 se
rect 2176 12104 2584 12376
tri 2584 12240 2720 12376 nw
tri 2720 12240 2856 12376 ne
tri 2584 12104 2720 12240 sw
tri 2720 12104 2856 12240 se
rect 2856 12104 3264 12376
tri 3264 12240 3400 12376 nw
tri 3264 12104 3400 12240 sw
rect 1360 11696 3400 12104
tri 1360 11560 1496 11696 ne
tri 1360 11424 1496 11560 se
rect 1496 11424 1904 11696
tri 1904 11560 2040 11696 nw
tri 2040 11560 2176 11696 ne
tri 1904 11424 2040 11560 sw
tri 2040 11424 2176 11560 se
rect 2176 11424 2584 11696
tri 2584 11560 2720 11696 nw
tri 2720 11560 2856 11696 ne
tri 2584 11424 2720 11560 sw
tri 2720 11424 2856 11560 se
rect 2856 11424 3264 11696
tri 3264 11560 3400 11696 nw
tri 3264 11424 3400 11560 sw
rect 1360 11016 3400 11424
tri 1360 10880 1496 11016 ne
rect 1496 10880 1904 11016
tri 1904 10880 2040 11016 nw
tri 2040 10880 2176 11016 ne
rect 2176 10880 2584 11016
tri 2584 10880 2720 11016 nw
tri 2720 10880 2856 11016 ne
rect 2856 10880 3264 11016
tri 3264 10880 3400 11016 nw
tri 4080 12784 4216 12920 se
rect 4216 12784 4624 13056
tri 4624 12920 4760 13056 nw
tri 6800 13464 6936 13600 se
rect 6936 13464 7344 13736
tri 7344 13600 7480 13736 nw
tri 8160 14144 8296 14280 se
rect 8296 14144 8704 14280
tri 8704 14144 8840 14280 sw
rect 8160 13736 8840 14144
tri 8160 13600 8296 13736 ne
rect 8296 13600 8704 13736
tri 8704 13600 8840 13736 nw
tri 9520 14144 9656 14280 se
rect 9656 14144 10064 14280
tri 10064 14144 10200 14280 sw
tri 10200 14144 10336 14280 se
rect 10336 14144 10744 14280
tri 10744 14144 10880 14280 sw
tri 10880 14144 11016 14280 se
rect 11016 14144 11424 14280
tri 11424 14144 11560 14280 sw
tri 11560 14144 11696 14280 se
rect 11696 14144 12104 14280
tri 12104 14144 12240 14280 sw
tri 12240 14144 12376 14280 se
rect 12376 14144 12784 14280
tri 12784 14144 12920 14280 sw
tri 12920 14144 13056 14280 se
rect 13056 14144 13464 14280
tri 13464 14144 13600 14280 sw
tri 13600 14144 13736 14280 se
rect 13736 14144 14144 14280
tri 14144 14144 14280 14280 sw
rect 9520 13736 14280 14144
tri 9520 13600 9656 13736 ne
tri 7344 13464 7480 13600 sw
tri 7480 13464 7616 13600 se
rect 7616 13464 8024 13600
tri 8024 13464 8160 13600 sw
rect 6800 13056 8160 13464
tri 6800 12920 6936 13056 ne
rect 6936 12920 7344 13056
tri 7344 12920 7480 13056 nw
tri 7480 12920 7616 13056 ne
tri 4624 12784 4760 12920 sw
rect 4080 12376 4760 12784
tri 4080 12240 4216 12376 ne
tri 4080 12104 4216 12240 se
rect 4216 12104 4624 12376
tri 4624 12240 4760 12376 nw
tri 7480 12784 7616 12920 se
rect 7616 12784 8024 13056
tri 8024 12920 8160 13056 nw
tri 9520 13464 9656 13600 se
rect 9656 13464 10064 13736
tri 10064 13600 10200 13736 nw
tri 10200 13600 10336 13736 ne
rect 10336 13600 10744 13736
tri 10744 13600 10880 13736 nw
tri 10880 13600 11016 13736 ne
rect 11016 13600 11424 13736
tri 11424 13600 11560 13736 nw
tri 11560 13600 11696 13736 ne
rect 11696 13600 12104 13736
tri 12104 13600 12240 13736 nw
tri 12240 13600 12376 13736 ne
rect 12376 13600 12784 13736
tri 12784 13600 12920 13736 nw
tri 12920 13600 13056 13736 ne
rect 13056 13600 13464 13736
tri 13464 13600 13600 13736 nw
tri 13600 13600 13736 13736 ne
tri 10064 13464 10200 13600 sw
rect 9520 13056 10200 13464
tri 9520 12920 9656 13056 ne
tri 8024 12784 8160 12920 sw
tri 8160 12784 8296 12920 se
rect 8296 12784 8704 12920
tri 8704 12784 8840 12920 sw
rect 7480 12376 8840 12784
tri 7480 12240 7616 12376 ne
tri 4624 12104 4760 12240 sw
rect 4080 11696 4760 12104
tri 4080 11560 4216 11696 ne
tri 4080 11424 4216 11560 se
rect 4216 11424 4624 11696
tri 4624 11560 4760 11696 nw
tri 6120 12104 6256 12240 se
rect 6256 12104 6664 12240
tri 6664 12104 6800 12240 sw
rect 6120 11696 6800 12104
tri 6120 11560 6256 11696 ne
tri 4624 11424 4760 11560 sw
rect 4080 11016 4760 11424
tri 4080 10880 4216 11016 ne
tri 544 10744 680 10880 sw
rect 0 10336 680 10744
tri 0 10200 136 10336 ne
tri 0 10064 136 10200 se
rect 136 10064 544 10336
tri 544 10200 680 10336 nw
tri 4080 10744 4216 10880 se
rect 4216 10744 4624 11016
tri 4624 10880 4760 11016 nw
tri 5440 11424 5576 11560 se
rect 5576 11424 5984 11560
tri 5984 11424 6120 11560 sw
tri 6120 11424 6256 11560 se
rect 6256 11424 6664 11696
tri 6664 11560 6800 11696 nw
tri 7480 12104 7616 12240 se
rect 7616 12104 8024 12376
tri 8024 12240 8160 12376 nw
tri 8160 12240 8296 12376 ne
tri 8024 12104 8160 12240 sw
tri 8160 12104 8296 12240 se
rect 8296 12104 8704 12376
tri 8704 12240 8840 12376 nw
tri 8704 12104 8840 12240 sw
rect 7480 11696 8840 12104
tri 7480 11560 7616 11696 ne
rect 7616 11560 8024 11696
tri 8024 11560 8160 11696 nw
tri 8160 11560 8296 11696 ne
rect 8296 11560 8704 11696
tri 8704 11560 8840 11696 nw
tri 9520 12784 9656 12920 se
rect 9656 12784 10064 13056
tri 10064 12920 10200 13056 nw
tri 13600 13464 13736 13600 se
rect 13736 13464 14144 13736
tri 14144 13600 14280 13736 nw
tri 14144 13464 14280 13600 sw
rect 13600 13056 14280 13464
tri 13600 12920 13736 13056 ne
tri 10064 12784 10200 12920 sw
rect 9520 12376 10200 12784
tri 9520 12240 9656 12376 ne
tri 9520 12104 9656 12240 se
rect 9656 12104 10064 12376
tri 10064 12240 10200 12376 nw
tri 10064 12104 10200 12240 sw
rect 9520 11696 10200 12104
tri 9520 11560 9656 11696 ne
tri 6664 11424 6800 11560 sw
rect 5440 11016 6800 11424
tri 5440 10880 5576 11016 ne
rect 5576 10880 5984 11016
tri 5984 10880 6120 11016 nw
tri 6120 10880 6256 11016 ne
tri 4624 10744 4760 10880 sw
rect 4080 10336 4760 10744
tri 4080 10200 4216 10336 ne
tri 544 10064 680 10200 sw
tri 680 10064 816 10200 se
rect 816 10064 1224 10200
tri 1224 10064 1360 10200 sw
tri 1360 10064 1496 10200 se
rect 1496 10064 1904 10200
tri 1904 10064 2040 10200 sw
tri 2040 10064 2176 10200 se
rect 2176 10064 2584 10200
tri 2584 10064 2720 10200 sw
tri 2720 10064 2856 10200 se
rect 2856 10064 3264 10200
tri 3264 10064 3400 10200 sw
tri 3400 10064 3536 10200 se
rect 3536 10064 3944 10200
tri 3944 10064 4080 10200 sw
tri 4080 10064 4216 10200 se
rect 4216 10064 4624 10336
tri 4624 10200 4760 10336 nw
tri 6120 10744 6256 10880 se
rect 6256 10744 6664 11016
tri 6664 10880 6800 11016 nw
tri 9520 11424 9656 11560 se
rect 9656 11424 10064 11696
tri 10064 11560 10200 11696 nw
tri 10064 11424 10200 11560 sw
rect 9520 11016 10200 11424
tri 9520 10880 9656 11016 ne
tri 6664 10744 6800 10880 sw
tri 6800 10744 6936 10880 se
rect 6936 10744 7344 10880
tri 7344 10744 7480 10880 sw
rect 6120 10336 7480 10744
tri 6120 10200 6256 10336 ne
rect 6256 10200 6664 10336
tri 6664 10200 6800 10336 nw
tri 6800 10200 6936 10336 ne
tri 4624 10064 4760 10200 sw
rect 0 9656 4760 10064
tri 0 9520 136 9656 ne
rect 136 9520 544 9656
tri 544 9520 680 9656 nw
tri 680 9520 816 9656 ne
rect 816 9520 1224 9656
tri 1224 9520 1360 9656 nw
tri 1360 9520 1496 9656 ne
rect 1496 9520 1904 9656
tri 1904 9520 2040 9656 nw
tri 2040 9520 2176 9656 ne
rect 2176 9520 2584 9656
tri 2584 9520 2720 9656 nw
tri 2720 9520 2856 9656 ne
rect 2856 9520 3264 9656
tri 3264 9520 3400 9656 nw
tri 3400 9520 3536 9656 ne
rect 3536 9520 3944 9656
tri 3944 9520 4080 9656 nw
tri 4080 9520 4216 9656 ne
rect 4216 9520 4624 9656
tri 4624 9520 4760 9656 nw
tri 5440 10064 5576 10200 se
rect 5576 10064 5984 10200
tri 5984 10064 6120 10200 sw
rect 5440 9656 6120 10064
tri 5440 9520 5576 9656 ne
tri 5440 9384 5576 9520 se
rect 5576 9384 5984 9656
tri 5984 9520 6120 9656 nw
tri 6800 10064 6936 10200 se
rect 6936 10064 7344 10336
tri 7344 10200 7480 10336 nw
tri 7344 10064 7480 10200 sw
rect 6800 9656 7480 10064
tri 6800 9520 6936 9656 ne
tri 5984 9384 6120 9520 sw
tri 6120 9384 6256 9520 se
rect 6256 9384 6664 9520
tri 6664 9384 6800 9520 sw
tri 6800 9384 6936 9520 se
rect 6936 9384 7344 9656
tri 7344 9520 7480 9656 nw
tri 8160 10744 8296 10880 se
rect 8296 10744 8704 10880
tri 8704 10744 8840 10880 sw
rect 8160 10336 8840 10744
tri 8160 10200 8296 10336 ne
tri 8160 10064 8296 10200 se
rect 8296 10064 8704 10336
tri 8704 10200 8840 10336 nw
tri 8704 10064 8840 10200 sw
rect 8160 9656 8840 10064
tri 8160 9520 8296 9656 ne
rect 8296 9520 8704 9656
tri 8704 9520 8840 9656 nw
tri 9520 10744 9656 10880 se
rect 9656 10744 10064 11016
tri 10064 10880 10200 11016 nw
tri 10880 12784 11016 12920 se
rect 11016 12784 11424 12920
tri 11424 12784 11560 12920 sw
tri 11560 12784 11696 12920 se
rect 11696 12784 12104 12920
tri 12104 12784 12240 12920 sw
tri 12240 12784 12376 12920 se
rect 12376 12784 12784 12920
tri 12784 12784 12920 12920 sw
rect 10880 12376 12920 12784
tri 10880 12240 11016 12376 ne
tri 10880 12104 11016 12240 se
rect 11016 12104 11424 12376
tri 11424 12240 11560 12376 nw
tri 11560 12240 11696 12376 ne
tri 11424 12104 11560 12240 sw
tri 11560 12104 11696 12240 se
rect 11696 12104 12104 12376
tri 12104 12240 12240 12376 nw
tri 12240 12240 12376 12376 ne
tri 12104 12104 12240 12240 sw
tri 12240 12104 12376 12240 se
rect 12376 12104 12784 12376
tri 12784 12240 12920 12376 nw
tri 12784 12104 12920 12240 sw
rect 10880 11696 12920 12104
tri 10880 11560 11016 11696 ne
tri 10880 11424 11016 11560 se
rect 11016 11424 11424 11696
tri 11424 11560 11560 11696 nw
tri 11560 11560 11696 11696 ne
tri 11424 11424 11560 11560 sw
tri 11560 11424 11696 11560 se
rect 11696 11424 12104 11696
tri 12104 11560 12240 11696 nw
tri 12240 11560 12376 11696 ne
tri 12104 11424 12240 11560 sw
tri 12240 11424 12376 11560 se
rect 12376 11424 12784 11696
tri 12784 11560 12920 11696 nw
tri 12784 11424 12920 11560 sw
rect 10880 11016 12920 11424
tri 10880 10880 11016 11016 ne
rect 11016 10880 11424 11016
tri 11424 10880 11560 11016 nw
tri 11560 10880 11696 11016 ne
rect 11696 10880 12104 11016
tri 12104 10880 12240 11016 nw
tri 12240 10880 12376 11016 ne
rect 12376 10880 12784 11016
tri 12784 10880 12920 11016 nw
tri 13600 12784 13736 12920 se
rect 13736 12784 14144 13056
tri 14144 12920 14280 13056 nw
tri 14144 12784 14280 12920 sw
rect 13600 12376 14280 12784
tri 13600 12240 13736 12376 ne
tri 13600 12104 13736 12240 se
rect 13736 12104 14144 12376
tri 14144 12240 14280 12376 nw
tri 14144 12104 14280 12240 sw
rect 13600 11696 14280 12104
tri 13600 11560 13736 11696 ne
tri 13600 11424 13736 11560 se
rect 13736 11424 14144 11696
tri 14144 11560 14280 11696 nw
tri 14144 11424 14280 11560 sw
rect 13600 11016 14280 11424
tri 13600 10880 13736 11016 ne
tri 10064 10744 10200 10880 sw
rect 9520 10336 10200 10744
tri 9520 10200 9656 10336 ne
tri 9520 10064 9656 10200 se
rect 9656 10064 10064 10336
tri 10064 10200 10200 10336 nw
tri 13600 10744 13736 10880 se
rect 13736 10744 14144 11016
tri 14144 10880 14280 11016 nw
tri 14144 10744 14280 10880 sw
rect 13600 10336 14280 10744
tri 13600 10200 13736 10336 ne
tri 10064 10064 10200 10200 sw
tri 10200 10064 10336 10200 se
rect 10336 10064 10744 10200
tri 10744 10064 10880 10200 sw
tri 10880 10064 11016 10200 se
rect 11016 10064 11424 10200
tri 11424 10064 11560 10200 sw
tri 11560 10064 11696 10200 se
rect 11696 10064 12104 10200
tri 12104 10064 12240 10200 sw
tri 12240 10064 12376 10200 se
rect 12376 10064 12784 10200
tri 12784 10064 12920 10200 sw
tri 12920 10064 13056 10200 se
rect 13056 10064 13464 10200
tri 13464 10064 13600 10200 sw
tri 13600 10064 13736 10200 se
rect 13736 10064 14144 10336
tri 14144 10200 14280 10336 nw
tri 14144 10064 14280 10200 sw
rect 9520 9656 14280 10064
tri 9520 9520 9656 9656 ne
rect 9656 9520 10064 9656
tri 10064 9520 10200 9656 nw
tri 10200 9520 10336 9656 ne
rect 10336 9520 10744 9656
tri 10744 9520 10880 9656 nw
tri 10880 9520 11016 9656 ne
rect 11016 9520 11424 9656
tri 11424 9520 11560 9656 nw
tri 11560 9520 11696 9656 ne
rect 11696 9520 12104 9656
tri 12104 9520 12240 9656 nw
tri 12240 9520 12376 9656 ne
rect 12376 9520 12784 9656
tri 12784 9520 12920 9656 nw
tri 12920 9520 13056 9656 ne
rect 13056 9520 13464 9656
tri 13464 9520 13600 9656 nw
tri 13600 9520 13736 9656 ne
rect 13736 9520 14144 9656
tri 14144 9520 14280 9656 nw
tri 7344 9384 7480 9520 sw
rect 5440 8976 7480 9384
tri 5440 8840 5576 8976 ne
tri 1360 8704 1496 8840 se
rect 1496 8704 1904 8840
tri 1904 8704 2040 8840 sw
tri 2040 8704 2176 8840 se
rect 2176 8704 2584 8840
tri 2584 8704 2720 8840 sw
rect 1360 8296 2720 8704
tri 1360 8160 1496 8296 ne
tri 1360 8024 1496 8160 se
rect 1496 8024 1904 8296
tri 1904 8160 2040 8296 nw
tri 2040 8160 2176 8296 ne
tri 1904 8024 2040 8160 sw
tri 2040 8024 2176 8160 se
rect 2176 8024 2584 8296
tri 2584 8160 2720 8296 nw
tri 4080 8704 4216 8840 se
rect 4216 8704 4624 8840
tri 4624 8704 4760 8840 sw
tri 4760 8704 4896 8840 se
rect 4896 8704 5304 8840
tri 5304 8704 5440 8840 sw
tri 5440 8704 5576 8840 se
rect 5576 8704 5984 8976
tri 5984 8840 6120 8976 nw
tri 6120 8840 6256 8976 ne
tri 5984 8704 6120 8840 sw
tri 6120 8704 6256 8840 se
rect 6256 8704 6664 8976
tri 6664 8840 6800 8976 nw
tri 6800 8840 6936 8976 ne
rect 6936 8840 7344 8976
tri 7344 8840 7480 8976 nw
tri 6664 8704 6800 8840 sw
rect 4080 8296 6800 8704
tri 4080 8160 4216 8296 ne
rect 4216 8160 4624 8296
tri 4624 8160 4760 8296 nw
tri 4760 8160 4896 8296 ne
tri 2584 8024 2720 8160 sw
rect 1360 7616 2720 8024
tri 1360 7480 1496 7616 ne
tri 0 7344 136 7480 se
rect 136 7344 544 7480
tri 544 7344 680 7480 sw
tri 680 7344 816 7480 se
rect 816 7344 1224 7480
tri 1224 7344 1360 7480 sw
tri 1360 7344 1496 7480 se
rect 1496 7344 1904 7616
tri 1904 7480 2040 7616 nw
tri 2040 7480 2176 7616 ne
tri 1904 7344 2040 7480 sw
tri 2040 7344 2176 7480 se
rect 2176 7344 2584 7616
tri 2584 7480 2720 7616 nw
tri 4760 8024 4896 8160 se
rect 4896 8024 5304 8296
tri 5304 8160 5440 8296 nw
tri 5440 8160 5576 8296 ne
tri 5304 8024 5440 8160 sw
tri 5440 8024 5576 8160 se
rect 5576 8024 5984 8296
tri 5984 8160 6120 8296 nw
tri 6120 8160 6256 8296 ne
tri 5984 8024 6120 8160 sw
tri 6120 8024 6256 8160 se
rect 6256 8024 6664 8296
tri 6664 8160 6800 8296 nw
tri 7480 8704 7616 8840 se
rect 7616 8704 8024 8840
tri 8024 8704 8160 8840 sw
rect 7480 8296 8160 8704
tri 7480 8160 7616 8296 ne
rect 7616 8160 8024 8296
tri 8024 8160 8160 8296 nw
tri 8840 8704 8976 8840 se
rect 8976 8704 9384 8840
tri 9384 8704 9520 8840 sw
tri 9520 8704 9656 8840 se
rect 9656 8704 10064 8840
tri 10064 8704 10200 8840 sw
rect 8840 8296 10200 8704
tri 8840 8160 8976 8296 ne
tri 6664 8024 6800 8160 sw
tri 6800 8024 6936 8160 se
rect 6936 8024 7344 8160
tri 7344 8024 7480 8160 sw
rect 4760 7616 7480 8024
tri 4760 7480 4896 7616 ne
tri 2584 7344 2720 7480 sw
tri 2720 7344 2856 7480 se
rect 2856 7344 3264 7480
tri 3264 7344 3400 7480 sw
tri 3400 7344 3536 7480 se
rect 3536 7344 3944 7480
tri 3944 7344 4080 7480 sw
tri 4080 7344 4216 7480 se
rect 4216 7344 4624 7480
tri 4624 7344 4760 7480 sw
tri 4760 7344 4896 7480 se
rect 4896 7344 5304 7616
tri 5304 7480 5440 7616 nw
tri 5440 7480 5576 7616 ne
rect 5576 7480 5984 7616
tri 5984 7480 6120 7616 nw
tri 6120 7480 6256 7616 ne
tri 5304 7344 5440 7480 sw
rect 0 6936 5440 7344
tri 0 6800 136 6936 ne
rect 136 6800 544 6936
tri 544 6800 680 6936 nw
tri 680 6800 816 6936 ne
tri 680 6664 816 6800 se
rect 816 6664 1224 6936
tri 1224 6800 1360 6936 nw
tri 1360 6800 1496 6936 ne
tri 1224 6664 1360 6800 sw
tri 1360 6664 1496 6800 se
rect 1496 6664 1904 6936
tri 1904 6800 2040 6936 nw
tri 2040 6800 2176 6936 ne
rect 2176 6800 2584 6936
tri 2584 6800 2720 6936 nw
tri 2720 6800 2856 6936 ne
tri 1904 6664 2040 6800 sw
rect 680 6256 2040 6664
tri 680 6120 816 6256 ne
rect 816 6120 1224 6256
tri 1224 6120 1360 6256 nw
tri 1360 6120 1496 6256 ne
rect 1496 6120 1904 6256
tri 1904 6120 2040 6256 nw
tri 2720 6664 2856 6800 se
rect 2856 6664 3264 6936
tri 3264 6800 3400 6936 nw
tri 3400 6800 3536 6936 ne
rect 3536 6800 3944 6936
tri 3944 6800 4080 6936 nw
tri 4080 6800 4216 6936 ne
rect 4216 6800 4624 6936
tri 4624 6800 4760 6936 nw
tri 4760 6800 4896 6936 ne
tri 3264 6664 3400 6800 sw
rect 2720 6256 3400 6664
tri 2720 6120 2856 6256 ne
tri 0 5984 136 6120 se
rect 136 5984 544 6120
tri 544 5984 680 6120 sw
rect 0 5576 680 5984
tri 0 5440 136 5576 ne
rect 136 5440 544 5576
tri 544 5440 680 5576 nw
tri 2720 5984 2856 6120 se
rect 2856 5984 3264 6256
tri 3264 6120 3400 6256 nw
tri 4760 6664 4896 6800 se
rect 4896 6664 5304 6936
tri 5304 6800 5440 6936 nw
tri 6120 7344 6256 7480 se
rect 6256 7344 6664 7616
tri 6664 7480 6800 7616 nw
tri 6800 7480 6936 7616 ne
rect 6936 7480 7344 7616
tri 7344 7480 7480 7616 nw
tri 8840 8024 8976 8160 se
rect 8976 8024 9384 8296
tri 9384 8160 9520 8296 nw
tri 9520 8160 9656 8296 ne
rect 9656 8160 10064 8296
tri 10064 8160 10200 8296 nw
tri 10880 8704 11016 8840 se
rect 11016 8704 11424 8840
tri 11424 8704 11560 8840 sw
rect 10880 8296 11560 8704
tri 10880 8160 11016 8296 ne
rect 11016 8160 11424 8296
tri 11424 8160 11560 8296 nw
tri 9384 8024 9520 8160 sw
rect 8840 7616 9520 8024
tri 8840 7480 8976 7616 ne
tri 6664 7344 6800 7480 sw
rect 6120 6936 6800 7344
tri 6120 6800 6256 6936 ne
tri 5304 6664 5440 6800 sw
tri 5440 6664 5576 6800 se
rect 5576 6664 5984 6800
tri 5984 6664 6120 6800 sw
tri 6120 6664 6256 6800 se
rect 6256 6664 6664 6936
tri 6664 6800 6800 6936 nw
tri 6664 6664 6800 6800 sw
rect 4760 6256 6800 6664
tri 4760 6120 4896 6256 ne
rect 4896 6120 5304 6256
tri 5304 6120 5440 6256 nw
tri 5440 6120 5576 6256 ne
tri 3264 5984 3400 6120 sw
tri 3400 5984 3536 6120 se
rect 3536 5984 3944 6120
tri 3944 5984 4080 6120 sw
tri 4080 5984 4216 6120 se
rect 4216 5984 4624 6120
tri 4624 5984 4760 6120 sw
rect 2720 5576 4760 5984
tri 2720 5440 2856 5576 ne
rect 2856 5440 3264 5576
tri 3264 5440 3400 5576 nw
tri 3400 5440 3536 5576 ne
rect 3536 5440 3944 5576
tri 3944 5440 4080 5576 nw
tri 4080 5440 4216 5576 ne
rect 4216 5440 4624 5576
tri 4624 5440 4760 5576 nw
tri 5440 5984 5576 6120 se
rect 5576 5984 5984 6256
tri 5984 6120 6120 6256 nw
tri 6120 6120 6256 6256 ne
tri 5984 5984 6120 6120 sw
tri 6120 5984 6256 6120 se
rect 6256 5984 6664 6256
tri 6664 6120 6800 6256 nw
tri 6664 5984 6800 6120 sw
rect 5440 5576 6800 5984
tri 5440 5440 5576 5576 ne
tri 5440 5304 5576 5440 se
rect 5576 5304 5984 5576
tri 5984 5440 6120 5576 nw
tri 6120 5440 6256 5576 ne
rect 6256 5440 6664 5576
tri 6664 5440 6800 5576 nw
tri 7480 7344 7616 7480 se
rect 7616 7344 8024 7480
tri 8024 7344 8160 7480 sw
rect 7480 6936 8160 7344
tri 7480 6800 7616 6936 ne
tri 7480 6664 7616 6800 se
rect 7616 6664 8024 6936
tri 8024 6800 8160 6936 nw
tri 8840 7344 8976 7480 se
rect 8976 7344 9384 7616
tri 9384 7480 9520 7616 nw
tri 9384 7344 9520 7480 sw
rect 8840 6936 9520 7344
tri 8840 6800 8976 6936 ne
tri 8024 6664 8160 6800 sw
tri 8160 6664 8296 6800 se
rect 8296 6664 8704 6800
tri 8704 6664 8840 6800 sw
tri 8840 6664 8976 6800 se
rect 8976 6664 9384 6936
tri 9384 6800 9520 6936 nw
tri 10200 8024 10336 8160 se
rect 10336 8024 10744 8160
tri 10744 8024 10880 8160 sw
rect 10200 7616 10880 8024
tri 10200 7480 10336 7616 ne
tri 10200 7344 10336 7480 se
rect 10336 7344 10744 7616
tri 10744 7480 10880 7616 nw
tri 12240 8024 12376 8160 se
rect 12376 8024 12784 8160
tri 12784 8024 12920 8160 sw
rect 12240 7616 12920 8024
tri 12240 7480 12376 7616 ne
rect 12376 7480 12784 7616
tri 12784 7480 12920 7616 nw
tri 10744 7344 10880 7480 sw
tri 10880 7344 11016 7480 se
rect 11016 7344 11424 7480
tri 11424 7344 11560 7480 sw
tri 11560 7344 11696 7480 se
rect 11696 7344 12104 7480
tri 12104 7344 12240 7480 sw
rect 10200 6936 12240 7344
tri 10200 6800 10336 6936 ne
rect 10336 6800 10744 6936
tri 10744 6800 10880 6936 nw
tri 10880 6800 11016 6936 ne
rect 11016 6800 11424 6936
tri 11424 6800 11560 6936 nw
tri 11560 6800 11696 6936 ne
rect 11696 6800 12104 6936
tri 12104 6800 12240 6936 nw
tri 13600 7344 13736 7480 se
rect 13736 7344 14144 7480
tri 14144 7344 14280 7480 sw
rect 13600 6936 14280 7344
tri 13600 6800 13736 6936 ne
rect 13736 6800 14144 6936
tri 14144 6800 14280 6936 nw
tri 9384 6664 9520 6800 sw
tri 9520 6664 9656 6800 se
rect 9656 6664 10064 6800
tri 10064 6664 10200 6800 sw
rect 7480 6256 10200 6664
tri 7480 6120 7616 6256 ne
tri 7480 5984 7616 6120 se
rect 7616 5984 8024 6256
tri 8024 6120 8160 6256 nw
tri 8160 6120 8296 6256 ne
tri 8024 5984 8160 6120 sw
tri 8160 5984 8296 6120 se
rect 8296 5984 8704 6256
tri 8704 6120 8840 6256 nw
tri 8840 6120 8976 6256 ne
rect 8976 6120 9384 6256
tri 9384 6120 9520 6256 nw
tri 9520 6120 9656 6256 ne
rect 9656 6120 10064 6256
tri 10064 6120 10200 6256 nw
tri 12920 6664 13056 6800 se
rect 13056 6664 13464 6800
tri 13464 6664 13600 6800 sw
rect 12920 6256 13600 6664
tri 12920 6120 13056 6256 ne
rect 13056 6120 13464 6256
tri 13464 6120 13600 6256 nw
tri 8704 5984 8840 6120 sw
rect 7480 5576 8840 5984
tri 7480 5440 7616 5576 ne
tri 5984 5304 6120 5440 sw
rect 5440 4896 6120 5304
tri 5440 4760 5576 4896 ne
tri 0 4624 136 4760 se
rect 136 4624 544 4760
tri 544 4624 680 4760 sw
tri 680 4624 816 4760 se
rect 816 4624 1224 4760
tri 1224 4624 1360 4760 sw
tri 1360 4624 1496 4760 se
rect 1496 4624 1904 4760
tri 1904 4624 2040 4760 sw
tri 2040 4624 2176 4760 se
rect 2176 4624 2584 4760
tri 2584 4624 2720 4760 sw
tri 2720 4624 2856 4760 se
rect 2856 4624 3264 4760
tri 3264 4624 3400 4760 sw
tri 3400 4624 3536 4760 se
rect 3536 4624 3944 4760
tri 3944 4624 4080 4760 sw
tri 4080 4624 4216 4760 se
rect 4216 4624 4624 4760
tri 4624 4624 4760 4760 sw
rect 0 4216 4760 4624
tri 0 4080 136 4216 ne
tri 0 3944 136 4080 se
rect 136 3944 544 4216
tri 544 4080 680 4216 nw
tri 680 4080 816 4216 ne
rect 816 4080 1224 4216
tri 1224 4080 1360 4216 nw
tri 1360 4080 1496 4216 ne
rect 1496 4080 1904 4216
tri 1904 4080 2040 4216 nw
tri 2040 4080 2176 4216 ne
rect 2176 4080 2584 4216
tri 2584 4080 2720 4216 nw
tri 2720 4080 2856 4216 ne
rect 2856 4080 3264 4216
tri 3264 4080 3400 4216 nw
tri 3400 4080 3536 4216 ne
rect 3536 4080 3944 4216
tri 3944 4080 4080 4216 nw
tri 4080 4080 4216 4216 ne
tri 544 3944 680 4080 sw
rect 0 3536 680 3944
tri 0 3400 136 3536 ne
tri 0 3264 136 3400 se
rect 136 3264 544 3536
tri 544 3400 680 3536 nw
tri 4080 3944 4216 4080 se
rect 4216 3944 4624 4216
tri 4624 4080 4760 4216 nw
tri 5440 4624 5576 4760 se
rect 5576 4624 5984 4896
tri 5984 4760 6120 4896 nw
tri 6800 5304 6936 5440 se
rect 6936 5304 7344 5440
tri 7344 5304 7480 5440 sw
tri 7480 5304 7616 5440 se
rect 7616 5304 8024 5576
tri 8024 5440 8160 5576 nw
tri 8160 5440 8296 5576 ne
tri 8024 5304 8160 5440 sw
tri 8160 5304 8296 5440 se
rect 8296 5304 8704 5576
tri 8704 5440 8840 5576 nw
tri 10880 5984 11016 6120 se
rect 11016 5984 11424 6120
tri 11424 5984 11560 6120 sw
rect 10880 5576 11560 5984
tri 10880 5440 11016 5576 ne
rect 11016 5440 11424 5576
tri 11424 5440 11560 5576 nw
tri 12240 5984 12376 6120 se
rect 12376 5984 12784 6120
tri 12784 5984 12920 6120 sw
rect 12240 5576 12920 5984
tri 12240 5440 12376 5576 ne
rect 12376 5440 12784 5576
tri 12784 5440 12920 5576 nw
tri 8704 5304 8840 5440 sw
tri 8840 5304 8976 5440 se
rect 8976 5304 9384 5440
tri 9384 5304 9520 5440 sw
rect 6800 4896 9520 5304
tri 6800 4760 6936 4896 ne
tri 5984 4624 6120 4760 sw
tri 6120 4624 6256 4760 se
rect 6256 4624 6664 4760
tri 6664 4624 6800 4760 sw
tri 6800 4624 6936 4760 se
rect 6936 4624 7344 4896
tri 7344 4760 7480 4896 nw
tri 7480 4760 7616 4896 ne
tri 7344 4624 7480 4760 sw
tri 7480 4624 7616 4760 se
rect 7616 4624 8024 4896
tri 8024 4760 8160 4896 nw
tri 8160 4760 8296 4896 ne
tri 8024 4624 8160 4760 sw
tri 8160 4624 8296 4760 se
rect 8296 4624 8704 4896
tri 8704 4760 8840 4896 nw
tri 8840 4760 8976 4896 ne
rect 8976 4760 9384 4896
tri 9384 4760 9520 4896 nw
tri 10200 5304 10336 5440 se
rect 10336 5304 10744 5440
tri 10744 5304 10880 5440 sw
rect 10200 4896 10880 5304
tri 10200 4760 10336 4896 ne
rect 10336 4760 10744 4896
tri 10744 4760 10880 4896 nw
tri 11560 5304 11696 5440 se
rect 11696 5304 12104 5440
tri 12104 5304 12240 5440 sw
rect 11560 4896 12240 5304
tri 11560 4760 11696 4896 ne
rect 11696 4760 12104 4896
tri 12104 4760 12240 4896 nw
tri 13600 5304 13736 5440 se
rect 13736 5304 14144 5440
tri 14144 5304 14280 5440 sw
rect 13600 4896 14280 5304
tri 13600 4760 13736 4896 ne
rect 13736 4760 14144 4896
tri 14144 4760 14280 4896 nw
tri 8704 4624 8840 4760 sw
rect 5440 4216 8840 4624
tri 5440 4080 5576 4216 ne
rect 5576 4080 5984 4216
tri 5984 4080 6120 4216 nw
tri 6120 4080 6256 4216 ne
rect 6256 4080 6664 4216
tri 6664 4080 6800 4216 nw
tri 6800 4080 6936 4216 ne
rect 6936 4080 7344 4216
tri 7344 4080 7480 4216 nw
tri 7480 4080 7616 4216 ne
rect 7616 4080 8024 4216
tri 8024 4080 8160 4216 nw
tri 8160 4080 8296 4216 ne
rect 8296 4080 8704 4216
tri 8704 4080 8840 4216 nw
tri 10880 4624 11016 4760 se
rect 11016 4624 11424 4760
tri 11424 4624 11560 4760 sw
rect 10880 4216 11560 4624
tri 10880 4080 11016 4216 ne
rect 11016 4080 11424 4216
tri 11424 4080 11560 4216 nw
tri 12920 4624 13056 4760 se
rect 13056 4624 13464 4760
tri 13464 4624 13600 4760 sw
rect 12920 4216 13600 4624
tri 12920 4080 13056 4216 ne
rect 13056 4080 13464 4216
tri 13464 4080 13600 4216 nw
tri 4624 3944 4760 4080 sw
rect 4080 3536 4760 3944
tri 4080 3400 4216 3536 ne
tri 544 3264 680 3400 sw
rect 0 2856 680 3264
tri 0 2720 136 2856 ne
tri 0 2584 136 2720 se
rect 136 2584 544 2856
tri 544 2720 680 2856 nw
tri 544 2584 680 2720 sw
rect 0 2176 680 2584
tri 0 2040 136 2176 ne
tri 0 1904 136 2040 se
rect 136 1904 544 2176
tri 544 2040 680 2176 nw
tri 544 1904 680 2040 sw
rect 0 1496 680 1904
tri 0 1360 136 1496 ne
tri 0 1224 136 1360 se
rect 136 1224 544 1496
tri 544 1360 680 1496 nw
tri 1360 3264 1496 3400 se
rect 1496 3264 1904 3400
tri 1904 3264 2040 3400 sw
tri 2040 3264 2176 3400 se
rect 2176 3264 2584 3400
tri 2584 3264 2720 3400 sw
tri 2720 3264 2856 3400 se
rect 2856 3264 3264 3400
tri 3264 3264 3400 3400 sw
rect 1360 2856 3400 3264
tri 1360 2720 1496 2856 ne
tri 1360 2584 1496 2720 se
rect 1496 2584 1904 2856
tri 1904 2720 2040 2856 nw
tri 2040 2720 2176 2856 ne
tri 1904 2584 2040 2720 sw
tri 2040 2584 2176 2720 se
rect 2176 2584 2584 2856
tri 2584 2720 2720 2856 nw
tri 2720 2720 2856 2856 ne
tri 2584 2584 2720 2720 sw
tri 2720 2584 2856 2720 se
rect 2856 2584 3264 2856
tri 3264 2720 3400 2856 nw
tri 3264 2584 3400 2720 sw
rect 1360 2176 3400 2584
tri 1360 2040 1496 2176 ne
tri 1360 1904 1496 2040 se
rect 1496 1904 1904 2176
tri 1904 2040 2040 2176 nw
tri 2040 2040 2176 2176 ne
tri 1904 1904 2040 2040 sw
tri 2040 1904 2176 2040 se
rect 2176 1904 2584 2176
tri 2584 2040 2720 2176 nw
tri 2720 2040 2856 2176 ne
tri 2584 1904 2720 2040 sw
tri 2720 1904 2856 2040 se
rect 2856 1904 3264 2176
tri 3264 2040 3400 2176 nw
tri 3264 1904 3400 2040 sw
rect 1360 1496 3400 1904
tri 1360 1360 1496 1496 ne
rect 1496 1360 1904 1496
tri 1904 1360 2040 1496 nw
tri 2040 1360 2176 1496 ne
rect 2176 1360 2584 1496
tri 2584 1360 2720 1496 nw
tri 2720 1360 2856 1496 ne
rect 2856 1360 3264 1496
tri 3264 1360 3400 1496 nw
tri 4080 3264 4216 3400 se
rect 4216 3264 4624 3536
tri 4624 3400 4760 3536 nw
tri 9520 3944 9656 4080 se
rect 9656 3944 10064 4080
tri 10064 3944 10200 4080 sw
rect 9520 3536 10200 3944
tri 9520 3400 9656 3536 ne
tri 4624 3264 4760 3400 sw
rect 4080 2856 4760 3264
tri 4080 2720 4216 2856 ne
tri 4080 2584 4216 2720 se
rect 4216 2584 4624 2856
tri 4624 2720 4760 2856 nw
tri 6120 3264 6256 3400 se
rect 6256 3264 6664 3400
tri 6664 3264 6800 3400 sw
tri 6800 3264 6936 3400 se
rect 6936 3264 7344 3400
tri 7344 3264 7480 3400 sw
tri 7480 3264 7616 3400 se
rect 7616 3264 8024 3400
tri 8024 3264 8160 3400 sw
rect 6120 2856 8160 3264
tri 6120 2720 6256 2856 ne
rect 6256 2720 6664 2856
tri 6664 2720 6800 2856 nw
tri 6800 2720 6936 2856 ne
tri 4624 2584 4760 2720 sw
rect 4080 2176 4760 2584
tri 4080 2040 4216 2176 ne
tri 4080 1904 4216 2040 se
rect 4216 1904 4624 2176
tri 4624 2040 4760 2176 nw
tri 4624 1904 4760 2040 sw
rect 4080 1496 4760 1904
tri 4080 1360 4216 1496 ne
tri 544 1224 680 1360 sw
rect 0 816 680 1224
tri 0 680 136 816 ne
tri 0 544 136 680 se
rect 136 544 544 816
tri 544 680 680 816 nw
tri 4080 1224 4216 1360 se
rect 4216 1224 4624 1496
tri 4624 1360 4760 1496 nw
tri 5440 2584 5576 2720 se
rect 5576 2584 5984 2720
tri 5984 2584 6120 2720 sw
rect 5440 2176 6120 2584
tri 5440 2040 5576 2176 ne
tri 5440 1904 5576 2040 se
rect 5576 1904 5984 2176
tri 5984 2040 6120 2176 nw
tri 6800 2584 6936 2720 se
rect 6936 2584 7344 2856
tri 7344 2720 7480 2856 nw
tri 7480 2720 7616 2856 ne
rect 7616 2720 8024 2856
tri 8024 2720 8160 2856 nw
tri 9520 3264 9656 3400 se
rect 9656 3264 10064 3536
tri 10064 3400 10200 3536 nw
tri 12240 3944 12376 4080 se
rect 12376 3944 12784 4080
tri 12784 3944 12920 4080 sw
rect 12240 3536 12920 3944
tri 12240 3400 12376 3536 ne
rect 12376 3400 12784 3536
tri 12784 3400 12920 3536 nw
tri 13600 3944 13736 4080 se
rect 13736 3944 14144 4080
tri 14144 3944 14280 4080 sw
rect 13600 3536 14280 3944
tri 13600 3400 13736 3536 ne
tri 10064 3264 10200 3400 sw
rect 9520 2856 10200 3264
tri 9520 2720 9656 2856 ne
tri 7344 2584 7480 2720 sw
rect 6800 2176 7480 2584
tri 6800 2040 6936 2176 ne
rect 6936 2040 7344 2176
tri 7344 2040 7480 2176 nw
tri 8160 2584 8296 2720 se
rect 8296 2584 8704 2720
tri 8704 2584 8840 2720 sw
rect 8160 2176 8840 2584
tri 8160 2040 8296 2176 ne
rect 8296 2040 8704 2176
tri 8704 2040 8840 2176 nw
tri 9520 2584 9656 2720 se
rect 9656 2584 10064 2856
tri 10064 2720 10200 2856 nw
tri 11560 3264 11696 3400 se
rect 11696 3264 12104 3400
tri 12104 3264 12240 3400 sw
rect 11560 2856 12240 3264
tri 11560 2720 11696 2856 ne
rect 11696 2720 12104 2856
tri 12104 2720 12240 2856 nw
tri 13600 3264 13736 3400 se
rect 13736 3264 14144 3536
tri 14144 3400 14280 3536 nw
tri 14144 3264 14280 3400 sw
rect 13600 2856 14280 3264
tri 13600 2720 13736 2856 ne
rect 13736 2720 14144 2856
tri 14144 2720 14280 2856 nw
tri 10064 2584 10200 2720 sw
rect 9520 2176 10200 2584
tri 9520 2040 9656 2176 ne
rect 9656 2040 10064 2176
tri 10064 2040 10200 2176 nw
tri 10880 2584 11016 2720 se
rect 11016 2584 11424 2720
tri 11424 2584 11560 2720 sw
rect 10880 2176 11560 2584
tri 10880 2040 11016 2176 ne
tri 5984 1904 6120 2040 sw
rect 5440 1496 6120 1904
tri 5440 1360 5576 1496 ne
rect 5576 1360 5984 1496
tri 5984 1360 6120 1496 nw
tri 7480 1904 7616 2040 se
rect 7616 1904 8024 2040
tri 8024 1904 8160 2040 sw
rect 7480 1496 8160 1904
tri 7480 1360 7616 1496 ne
tri 4624 1224 4760 1360 sw
rect 4080 816 4760 1224
tri 4080 680 4216 816 ne
tri 544 544 680 680 sw
tri 680 544 816 680 se
rect 816 544 1224 680
tri 1224 544 1360 680 sw
tri 1360 544 1496 680 se
rect 1496 544 1904 680
tri 1904 544 2040 680 sw
tri 2040 544 2176 680 se
rect 2176 544 2584 680
tri 2584 544 2720 680 sw
tri 2720 544 2856 680 se
rect 2856 544 3264 680
tri 3264 544 3400 680 sw
tri 3400 544 3536 680 se
rect 3536 544 3944 680
tri 3944 544 4080 680 sw
tri 4080 544 4216 680 se
rect 4216 544 4624 816
tri 4624 680 4760 816 nw
tri 6120 1224 6256 1360 se
rect 6256 1224 6664 1360
tri 6664 1224 6800 1360 sw
tri 6800 1224 6936 1360 se
rect 6936 1224 7344 1360
tri 7344 1224 7480 1360 sw
tri 7480 1224 7616 1360 se
rect 7616 1224 8024 1496
tri 8024 1360 8160 1496 nw
tri 10880 1904 11016 2040 se
rect 11016 1904 11424 2176
tri 11424 2040 11560 2176 nw
tri 12920 2584 13056 2720 se
rect 13056 2584 13464 2720
tri 13464 2584 13600 2720 sw
rect 12920 2176 13600 2584
tri 12920 2040 13056 2176 ne
rect 13056 2040 13464 2176
tri 13464 2040 13600 2176 nw
tri 11424 1904 11560 2040 sw
rect 10880 1496 11560 1904
tri 10880 1360 11016 1496 ne
tri 8024 1224 8160 1360 sw
rect 6120 816 8160 1224
tri 6120 680 6256 816 ne
rect 6256 680 6664 816
tri 6664 680 6800 816 nw
tri 6800 680 6936 816 ne
rect 6936 680 7344 816
tri 7344 680 7480 816 nw
tri 7480 680 7616 816 ne
rect 7616 680 8024 816
tri 8024 680 8160 816 nw
tri 8840 1224 8976 1360 se
rect 8976 1224 9384 1360
tri 9384 1224 9520 1360 sw
rect 8840 816 9520 1224
tri 8840 680 8976 816 ne
rect 8976 680 9384 816
tri 9384 680 9520 816 nw
tri 10880 1224 11016 1360 se
rect 11016 1224 11424 1496
tri 11424 1360 11560 1496 nw
tri 12240 1904 12376 2040 se
rect 12376 1904 12784 2040
tri 12784 1904 12920 2040 sw
rect 12240 1496 12920 1904
tri 12240 1360 12376 1496 ne
rect 12376 1360 12784 1496
tri 12784 1360 12920 1496 nw
tri 11424 1224 11560 1360 sw
tri 11560 1224 11696 1360 se
rect 11696 1224 12104 1360
tri 12104 1224 12240 1360 sw
rect 10880 816 12240 1224
tri 10880 680 11016 816 ne
rect 11016 680 11424 816
tri 11424 680 11560 816 nw
tri 11560 680 11696 816 ne
rect 11696 680 12104 816
tri 12104 680 12240 816 nw
tri 12920 1224 13056 1360 se
rect 13056 1224 13464 1360
tri 13464 1224 13600 1360 sw
tri 13600 1224 13736 1360 se
rect 13736 1224 14144 1360
tri 14144 1224 14280 1360 sw
rect 12920 816 14280 1224
tri 12920 680 13056 816 ne
tri 4624 544 4760 680 sw
rect 0 136 4760 544
tri 0 0 136 136 ne
rect 136 0 544 136
tri 544 0 680 136 nw
tri 680 0 816 136 ne
rect 816 0 1224 136
tri 1224 0 1360 136 nw
tri 1360 0 1496 136 ne
rect 1496 0 1904 136
tri 1904 0 2040 136 nw
tri 2040 0 2176 136 ne
rect 2176 0 2584 136
tri 2584 0 2720 136 nw
tri 2720 0 2856 136 ne
rect 2856 0 3264 136
tri 3264 0 3400 136 nw
tri 3400 0 3536 136 ne
rect 3536 0 3944 136
tri 3944 0 4080 136 nw
tri 4080 0 4216 136 ne
rect 4216 0 4624 136
tri 4624 0 4760 136 nw
tri 8160 544 8296 680 se
rect 8296 544 8704 680
tri 8704 544 8840 680 sw
rect 8160 136 8840 544
tri 8160 0 8296 136 ne
rect 8296 0 8704 136
tri 8704 0 8840 136 nw
tri 10200 544 10336 680 se
rect 10336 544 10744 680
tri 10744 544 10880 680 sw
rect 10200 136 10880 544
tri 10200 0 10336 136 ne
rect 10336 0 10744 136
tri 10744 0 10880 136 nw
tri 12920 544 13056 680 se
rect 13056 544 13464 816
tri 13464 680 13600 816 nw
tri 13600 680 13736 816 ne
rect 13736 680 14144 816
tri 14144 680 14280 816 nw
tri 13464 544 13600 680 sw
rect 12920 136 13600 544
tri 12920 0 13056 136 ne
rect 13056 0 13464 136
tri 13464 0 13600 136 nw
<< metal3 >>
tri 0 14144 136 14280 se
rect 136 14144 544 14280
tri 544 14144 680 14280 sw
tri 680 14144 816 14280 se
rect 816 14144 1224 14280
tri 1224 14144 1360 14280 sw
tri 1360 14144 1496 14280 se
rect 1496 14144 1904 14280
tri 1904 14144 2040 14280 sw
tri 2040 14144 2176 14280 se
rect 2176 14144 2584 14280
tri 2584 14144 2720 14280 sw
tri 2720 14144 2856 14280 se
rect 2856 14144 3264 14280
tri 3264 14144 3400 14280 sw
tri 3400 14144 3536 14280 se
rect 3536 14144 3944 14280
tri 3944 14144 4080 14280 sw
tri 4080 14144 4216 14280 se
rect 4216 14144 4624 14280
tri 4624 14144 4760 14280 sw
rect 0 13736 4760 14144
tri 0 13600 136 13736 ne
tri 0 13464 136 13600 se
rect 136 13464 544 13736
tri 544 13600 680 13736 nw
tri 680 13600 816 13736 ne
rect 816 13600 1224 13736
tri 1224 13600 1360 13736 nw
tri 1360 13600 1496 13736 ne
rect 1496 13600 1904 13736
tri 1904 13600 2040 13736 nw
tri 2040 13600 2176 13736 ne
rect 2176 13600 2584 13736
tri 2584 13600 2720 13736 nw
tri 2720 13600 2856 13736 ne
rect 2856 13600 3264 13736
tri 3264 13600 3400 13736 nw
tri 3400 13600 3536 13736 ne
rect 3536 13600 3944 13736
tri 3944 13600 4080 13736 nw
tri 4080 13600 4216 13736 ne
tri 544 13464 680 13600 sw
rect 0 13056 680 13464
tri 0 12920 136 13056 ne
tri 0 12784 136 12920 se
rect 136 12784 544 13056
tri 544 12920 680 13056 nw
tri 4080 13464 4216 13600 se
rect 4216 13464 4624 13736
tri 4624 13600 4760 13736 nw
tri 6120 14144 6256 14280 se
rect 6256 14144 6664 14280
tri 6664 14144 6800 14280 sw
tri 6800 14144 6936 14280 se
rect 6936 14144 7344 14280
tri 7344 14144 7480 14280 sw
rect 6120 13736 7480 14144
tri 6120 13600 6256 13736 ne
rect 6256 13600 6664 13736
tri 6664 13600 6800 13736 nw
tri 6800 13600 6936 13736 ne
tri 4624 13464 4760 13600 sw
rect 4080 13056 4760 13464
tri 4080 12920 4216 13056 ne
tri 544 12784 680 12920 sw
rect 0 12376 680 12784
tri 0 12240 136 12376 ne
tri 0 12104 136 12240 se
rect 136 12104 544 12376
tri 544 12240 680 12376 nw
tri 544 12104 680 12240 sw
rect 0 11696 680 12104
tri 0 11560 136 11696 ne
tri 0 11424 136 11560 se
rect 136 11424 544 11696
tri 544 11560 680 11696 nw
tri 544 11424 680 11560 sw
rect 0 11016 680 11424
tri 0 10880 136 11016 ne
tri 0 10744 136 10880 se
rect 136 10744 544 11016
tri 544 10880 680 11016 nw
tri 1360 12784 1496 12920 se
rect 1496 12784 1904 12920
tri 1904 12784 2040 12920 sw
tri 2040 12784 2176 12920 se
rect 2176 12784 2584 12920
tri 2584 12784 2720 12920 sw
tri 2720 12784 2856 12920 se
rect 2856 12784 3264 12920
tri 3264 12784 3400 12920 sw
rect 1360 12376 3400 12784
tri 1360 12240 1496 12376 ne
tri 1360 12104 1496 12240 se
rect 1496 12104 1904 12376
tri 1904 12240 2040 12376 nw
tri 2040 12240 2176 12376 ne
tri 1904 12104 2040 12240 sw
tri 2040 12104 2176 12240 se
rect 2176 12104 2584 12376
tri 2584 12240 2720 12376 nw
tri 2720 12240 2856 12376 ne
tri 2584 12104 2720 12240 sw
tri 2720 12104 2856 12240 se
rect 2856 12104 3264 12376
tri 3264 12240 3400 12376 nw
tri 3264 12104 3400 12240 sw
rect 1360 11696 3400 12104
tri 1360 11560 1496 11696 ne
tri 1360 11424 1496 11560 se
rect 1496 11424 1904 11696
tri 1904 11560 2040 11696 nw
tri 2040 11560 2176 11696 ne
tri 1904 11424 2040 11560 sw
tri 2040 11424 2176 11560 se
rect 2176 11424 2584 11696
tri 2584 11560 2720 11696 nw
tri 2720 11560 2856 11696 ne
tri 2584 11424 2720 11560 sw
tri 2720 11424 2856 11560 se
rect 2856 11424 3264 11696
tri 3264 11560 3400 11696 nw
tri 3264 11424 3400 11560 sw
rect 1360 11016 3400 11424
tri 1360 10880 1496 11016 ne
rect 1496 10880 1904 11016
tri 1904 10880 2040 11016 nw
tri 2040 10880 2176 11016 ne
rect 2176 10880 2584 11016
tri 2584 10880 2720 11016 nw
tri 2720 10880 2856 11016 ne
rect 2856 10880 3264 11016
tri 3264 10880 3400 11016 nw
tri 4080 12784 4216 12920 se
rect 4216 12784 4624 13056
tri 4624 12920 4760 13056 nw
tri 6800 13464 6936 13600 se
rect 6936 13464 7344 13736
tri 7344 13600 7480 13736 nw
tri 8160 14144 8296 14280 se
rect 8296 14144 8704 14280
tri 8704 14144 8840 14280 sw
rect 8160 13736 8840 14144
tri 8160 13600 8296 13736 ne
rect 8296 13600 8704 13736
tri 8704 13600 8840 13736 nw
tri 9520 14144 9656 14280 se
rect 9656 14144 10064 14280
tri 10064 14144 10200 14280 sw
tri 10200 14144 10336 14280 se
rect 10336 14144 10744 14280
tri 10744 14144 10880 14280 sw
tri 10880 14144 11016 14280 se
rect 11016 14144 11424 14280
tri 11424 14144 11560 14280 sw
tri 11560 14144 11696 14280 se
rect 11696 14144 12104 14280
tri 12104 14144 12240 14280 sw
tri 12240 14144 12376 14280 se
rect 12376 14144 12784 14280
tri 12784 14144 12920 14280 sw
tri 12920 14144 13056 14280 se
rect 13056 14144 13464 14280
tri 13464 14144 13600 14280 sw
tri 13600 14144 13736 14280 se
rect 13736 14144 14144 14280
tri 14144 14144 14280 14280 sw
rect 9520 13736 14280 14144
tri 9520 13600 9656 13736 ne
tri 7344 13464 7480 13600 sw
tri 7480 13464 7616 13600 se
rect 7616 13464 8024 13600
tri 8024 13464 8160 13600 sw
rect 6800 13056 8160 13464
tri 6800 12920 6936 13056 ne
rect 6936 12920 7344 13056
tri 7344 12920 7480 13056 nw
tri 7480 12920 7616 13056 ne
tri 4624 12784 4760 12920 sw
rect 4080 12376 4760 12784
tri 4080 12240 4216 12376 ne
tri 4080 12104 4216 12240 se
rect 4216 12104 4624 12376
tri 4624 12240 4760 12376 nw
tri 7480 12784 7616 12920 se
rect 7616 12784 8024 13056
tri 8024 12920 8160 13056 nw
tri 9520 13464 9656 13600 se
rect 9656 13464 10064 13736
tri 10064 13600 10200 13736 nw
tri 10200 13600 10336 13736 ne
rect 10336 13600 10744 13736
tri 10744 13600 10880 13736 nw
tri 10880 13600 11016 13736 ne
rect 11016 13600 11424 13736
tri 11424 13600 11560 13736 nw
tri 11560 13600 11696 13736 ne
rect 11696 13600 12104 13736
tri 12104 13600 12240 13736 nw
tri 12240 13600 12376 13736 ne
rect 12376 13600 12784 13736
tri 12784 13600 12920 13736 nw
tri 12920 13600 13056 13736 ne
rect 13056 13600 13464 13736
tri 13464 13600 13600 13736 nw
tri 13600 13600 13736 13736 ne
tri 10064 13464 10200 13600 sw
rect 9520 13056 10200 13464
tri 9520 12920 9656 13056 ne
tri 8024 12784 8160 12920 sw
tri 8160 12784 8296 12920 se
rect 8296 12784 8704 12920
tri 8704 12784 8840 12920 sw
rect 7480 12376 8840 12784
tri 7480 12240 7616 12376 ne
tri 4624 12104 4760 12240 sw
rect 4080 11696 4760 12104
tri 4080 11560 4216 11696 ne
tri 4080 11424 4216 11560 se
rect 4216 11424 4624 11696
tri 4624 11560 4760 11696 nw
tri 6120 12104 6256 12240 se
rect 6256 12104 6664 12240
tri 6664 12104 6800 12240 sw
rect 6120 11696 6800 12104
tri 6120 11560 6256 11696 ne
tri 4624 11424 4760 11560 sw
rect 4080 11016 4760 11424
tri 4080 10880 4216 11016 ne
tri 544 10744 680 10880 sw
rect 0 10336 680 10744
tri 0 10200 136 10336 ne
tri 0 10064 136 10200 se
rect 136 10064 544 10336
tri 544 10200 680 10336 nw
tri 4080 10744 4216 10880 se
rect 4216 10744 4624 11016
tri 4624 10880 4760 11016 nw
tri 5440 11424 5576 11560 se
rect 5576 11424 5984 11560
tri 5984 11424 6120 11560 sw
tri 6120 11424 6256 11560 se
rect 6256 11424 6664 11696
tri 6664 11560 6800 11696 nw
tri 7480 12104 7616 12240 se
rect 7616 12104 8024 12376
tri 8024 12240 8160 12376 nw
tri 8160 12240 8296 12376 ne
tri 8024 12104 8160 12240 sw
tri 8160 12104 8296 12240 se
rect 8296 12104 8704 12376
tri 8704 12240 8840 12376 nw
tri 8704 12104 8840 12240 sw
rect 7480 11696 8840 12104
tri 7480 11560 7616 11696 ne
rect 7616 11560 8024 11696
tri 8024 11560 8160 11696 nw
tri 8160 11560 8296 11696 ne
rect 8296 11560 8704 11696
tri 8704 11560 8840 11696 nw
tri 9520 12784 9656 12920 se
rect 9656 12784 10064 13056
tri 10064 12920 10200 13056 nw
tri 13600 13464 13736 13600 se
rect 13736 13464 14144 13736
tri 14144 13600 14280 13736 nw
tri 14144 13464 14280 13600 sw
rect 13600 13056 14280 13464
tri 13600 12920 13736 13056 ne
tri 10064 12784 10200 12920 sw
rect 9520 12376 10200 12784
tri 9520 12240 9656 12376 ne
tri 9520 12104 9656 12240 se
rect 9656 12104 10064 12376
tri 10064 12240 10200 12376 nw
tri 10064 12104 10200 12240 sw
rect 9520 11696 10200 12104
tri 9520 11560 9656 11696 ne
tri 6664 11424 6800 11560 sw
rect 5440 11016 6800 11424
tri 5440 10880 5576 11016 ne
rect 5576 10880 5984 11016
tri 5984 10880 6120 11016 nw
tri 6120 10880 6256 11016 ne
tri 4624 10744 4760 10880 sw
rect 4080 10336 4760 10744
tri 4080 10200 4216 10336 ne
tri 544 10064 680 10200 sw
tri 680 10064 816 10200 se
rect 816 10064 1224 10200
tri 1224 10064 1360 10200 sw
tri 1360 10064 1496 10200 se
rect 1496 10064 1904 10200
tri 1904 10064 2040 10200 sw
tri 2040 10064 2176 10200 se
rect 2176 10064 2584 10200
tri 2584 10064 2720 10200 sw
tri 2720 10064 2856 10200 se
rect 2856 10064 3264 10200
tri 3264 10064 3400 10200 sw
tri 3400 10064 3536 10200 se
rect 3536 10064 3944 10200
tri 3944 10064 4080 10200 sw
tri 4080 10064 4216 10200 se
rect 4216 10064 4624 10336
tri 4624 10200 4760 10336 nw
tri 6120 10744 6256 10880 se
rect 6256 10744 6664 11016
tri 6664 10880 6800 11016 nw
tri 9520 11424 9656 11560 se
rect 9656 11424 10064 11696
tri 10064 11560 10200 11696 nw
tri 10064 11424 10200 11560 sw
rect 9520 11016 10200 11424
tri 9520 10880 9656 11016 ne
tri 6664 10744 6800 10880 sw
tri 6800 10744 6936 10880 se
rect 6936 10744 7344 10880
tri 7344 10744 7480 10880 sw
rect 6120 10336 7480 10744
tri 6120 10200 6256 10336 ne
rect 6256 10200 6664 10336
tri 6664 10200 6800 10336 nw
tri 6800 10200 6936 10336 ne
tri 4624 10064 4760 10200 sw
rect 0 9656 4760 10064
tri 0 9520 136 9656 ne
rect 136 9520 544 9656
tri 544 9520 680 9656 nw
tri 680 9520 816 9656 ne
rect 816 9520 1224 9656
tri 1224 9520 1360 9656 nw
tri 1360 9520 1496 9656 ne
rect 1496 9520 1904 9656
tri 1904 9520 2040 9656 nw
tri 2040 9520 2176 9656 ne
rect 2176 9520 2584 9656
tri 2584 9520 2720 9656 nw
tri 2720 9520 2856 9656 ne
rect 2856 9520 3264 9656
tri 3264 9520 3400 9656 nw
tri 3400 9520 3536 9656 ne
rect 3536 9520 3944 9656
tri 3944 9520 4080 9656 nw
tri 4080 9520 4216 9656 ne
rect 4216 9520 4624 9656
tri 4624 9520 4760 9656 nw
tri 5440 10064 5576 10200 se
rect 5576 10064 5984 10200
tri 5984 10064 6120 10200 sw
rect 5440 9656 6120 10064
tri 5440 9520 5576 9656 ne
tri 5440 9384 5576 9520 se
rect 5576 9384 5984 9656
tri 5984 9520 6120 9656 nw
tri 6800 10064 6936 10200 se
rect 6936 10064 7344 10336
tri 7344 10200 7480 10336 nw
tri 7344 10064 7480 10200 sw
rect 6800 9656 7480 10064
tri 6800 9520 6936 9656 ne
tri 5984 9384 6120 9520 sw
tri 6120 9384 6256 9520 se
rect 6256 9384 6664 9520
tri 6664 9384 6800 9520 sw
tri 6800 9384 6936 9520 se
rect 6936 9384 7344 9656
tri 7344 9520 7480 9656 nw
tri 8160 10744 8296 10880 se
rect 8296 10744 8704 10880
tri 8704 10744 8840 10880 sw
rect 8160 10336 8840 10744
tri 8160 10200 8296 10336 ne
tri 8160 10064 8296 10200 se
rect 8296 10064 8704 10336
tri 8704 10200 8840 10336 nw
tri 8704 10064 8840 10200 sw
rect 8160 9656 8840 10064
tri 8160 9520 8296 9656 ne
rect 8296 9520 8704 9656
tri 8704 9520 8840 9656 nw
tri 9520 10744 9656 10880 se
rect 9656 10744 10064 11016
tri 10064 10880 10200 11016 nw
tri 10880 12784 11016 12920 se
rect 11016 12784 11424 12920
tri 11424 12784 11560 12920 sw
tri 11560 12784 11696 12920 se
rect 11696 12784 12104 12920
tri 12104 12784 12240 12920 sw
tri 12240 12784 12376 12920 se
rect 12376 12784 12784 12920
tri 12784 12784 12920 12920 sw
rect 10880 12376 12920 12784
tri 10880 12240 11016 12376 ne
tri 10880 12104 11016 12240 se
rect 11016 12104 11424 12376
tri 11424 12240 11560 12376 nw
tri 11560 12240 11696 12376 ne
tri 11424 12104 11560 12240 sw
tri 11560 12104 11696 12240 se
rect 11696 12104 12104 12376
tri 12104 12240 12240 12376 nw
tri 12240 12240 12376 12376 ne
tri 12104 12104 12240 12240 sw
tri 12240 12104 12376 12240 se
rect 12376 12104 12784 12376
tri 12784 12240 12920 12376 nw
tri 12784 12104 12920 12240 sw
rect 10880 11696 12920 12104
tri 10880 11560 11016 11696 ne
tri 10880 11424 11016 11560 se
rect 11016 11424 11424 11696
tri 11424 11560 11560 11696 nw
tri 11560 11560 11696 11696 ne
tri 11424 11424 11560 11560 sw
tri 11560 11424 11696 11560 se
rect 11696 11424 12104 11696
tri 12104 11560 12240 11696 nw
tri 12240 11560 12376 11696 ne
tri 12104 11424 12240 11560 sw
tri 12240 11424 12376 11560 se
rect 12376 11424 12784 11696
tri 12784 11560 12920 11696 nw
tri 12784 11424 12920 11560 sw
rect 10880 11016 12920 11424
tri 10880 10880 11016 11016 ne
rect 11016 10880 11424 11016
tri 11424 10880 11560 11016 nw
tri 11560 10880 11696 11016 ne
rect 11696 10880 12104 11016
tri 12104 10880 12240 11016 nw
tri 12240 10880 12376 11016 ne
rect 12376 10880 12784 11016
tri 12784 10880 12920 11016 nw
tri 13600 12784 13736 12920 se
rect 13736 12784 14144 13056
tri 14144 12920 14280 13056 nw
tri 14144 12784 14280 12920 sw
rect 13600 12376 14280 12784
tri 13600 12240 13736 12376 ne
tri 13600 12104 13736 12240 se
rect 13736 12104 14144 12376
tri 14144 12240 14280 12376 nw
tri 14144 12104 14280 12240 sw
rect 13600 11696 14280 12104
tri 13600 11560 13736 11696 ne
tri 13600 11424 13736 11560 se
rect 13736 11424 14144 11696
tri 14144 11560 14280 11696 nw
tri 14144 11424 14280 11560 sw
rect 13600 11016 14280 11424
tri 13600 10880 13736 11016 ne
tri 10064 10744 10200 10880 sw
rect 9520 10336 10200 10744
tri 9520 10200 9656 10336 ne
tri 9520 10064 9656 10200 se
rect 9656 10064 10064 10336
tri 10064 10200 10200 10336 nw
tri 13600 10744 13736 10880 se
rect 13736 10744 14144 11016
tri 14144 10880 14280 11016 nw
tri 14144 10744 14280 10880 sw
rect 13600 10336 14280 10744
tri 13600 10200 13736 10336 ne
tri 10064 10064 10200 10200 sw
tri 10200 10064 10336 10200 se
rect 10336 10064 10744 10200
tri 10744 10064 10880 10200 sw
tri 10880 10064 11016 10200 se
rect 11016 10064 11424 10200
tri 11424 10064 11560 10200 sw
tri 11560 10064 11696 10200 se
rect 11696 10064 12104 10200
tri 12104 10064 12240 10200 sw
tri 12240 10064 12376 10200 se
rect 12376 10064 12784 10200
tri 12784 10064 12920 10200 sw
tri 12920 10064 13056 10200 se
rect 13056 10064 13464 10200
tri 13464 10064 13600 10200 sw
tri 13600 10064 13736 10200 se
rect 13736 10064 14144 10336
tri 14144 10200 14280 10336 nw
tri 14144 10064 14280 10200 sw
rect 9520 9656 14280 10064
tri 9520 9520 9656 9656 ne
rect 9656 9520 10064 9656
tri 10064 9520 10200 9656 nw
tri 10200 9520 10336 9656 ne
rect 10336 9520 10744 9656
tri 10744 9520 10880 9656 nw
tri 10880 9520 11016 9656 ne
rect 11016 9520 11424 9656
tri 11424 9520 11560 9656 nw
tri 11560 9520 11696 9656 ne
rect 11696 9520 12104 9656
tri 12104 9520 12240 9656 nw
tri 12240 9520 12376 9656 ne
rect 12376 9520 12784 9656
tri 12784 9520 12920 9656 nw
tri 12920 9520 13056 9656 ne
rect 13056 9520 13464 9656
tri 13464 9520 13600 9656 nw
tri 13600 9520 13736 9656 ne
rect 13736 9520 14144 9656
tri 14144 9520 14280 9656 nw
tri 7344 9384 7480 9520 sw
rect 5440 8976 7480 9384
tri 5440 8840 5576 8976 ne
tri 1360 8704 1496 8840 se
rect 1496 8704 1904 8840
tri 1904 8704 2040 8840 sw
tri 2040 8704 2176 8840 se
rect 2176 8704 2584 8840
tri 2584 8704 2720 8840 sw
rect 1360 8296 2720 8704
tri 1360 8160 1496 8296 ne
tri 1360 8024 1496 8160 se
rect 1496 8024 1904 8296
tri 1904 8160 2040 8296 nw
tri 2040 8160 2176 8296 ne
tri 1904 8024 2040 8160 sw
tri 2040 8024 2176 8160 se
rect 2176 8024 2584 8296
tri 2584 8160 2720 8296 nw
tri 4080 8704 4216 8840 se
rect 4216 8704 4624 8840
tri 4624 8704 4760 8840 sw
tri 4760 8704 4896 8840 se
rect 4896 8704 5304 8840
tri 5304 8704 5440 8840 sw
tri 5440 8704 5576 8840 se
rect 5576 8704 5984 8976
tri 5984 8840 6120 8976 nw
tri 6120 8840 6256 8976 ne
tri 5984 8704 6120 8840 sw
tri 6120 8704 6256 8840 se
rect 6256 8704 6664 8976
tri 6664 8840 6800 8976 nw
tri 6800 8840 6936 8976 ne
rect 6936 8840 7344 8976
tri 7344 8840 7480 8976 nw
tri 6664 8704 6800 8840 sw
rect 4080 8296 6800 8704
tri 4080 8160 4216 8296 ne
rect 4216 8160 4624 8296
tri 4624 8160 4760 8296 nw
tri 4760 8160 4896 8296 ne
tri 2584 8024 2720 8160 sw
rect 1360 7616 2720 8024
tri 1360 7480 1496 7616 ne
tri 0 7344 136 7480 se
rect 136 7344 544 7480
tri 544 7344 680 7480 sw
tri 680 7344 816 7480 se
rect 816 7344 1224 7480
tri 1224 7344 1360 7480 sw
tri 1360 7344 1496 7480 se
rect 1496 7344 1904 7616
tri 1904 7480 2040 7616 nw
tri 2040 7480 2176 7616 ne
tri 1904 7344 2040 7480 sw
tri 2040 7344 2176 7480 se
rect 2176 7344 2584 7616
tri 2584 7480 2720 7616 nw
tri 4760 8024 4896 8160 se
rect 4896 8024 5304 8296
tri 5304 8160 5440 8296 nw
tri 5440 8160 5576 8296 ne
tri 5304 8024 5440 8160 sw
tri 5440 8024 5576 8160 se
rect 5576 8024 5984 8296
tri 5984 8160 6120 8296 nw
tri 6120 8160 6256 8296 ne
tri 5984 8024 6120 8160 sw
tri 6120 8024 6256 8160 se
rect 6256 8024 6664 8296
tri 6664 8160 6800 8296 nw
tri 7480 8704 7616 8840 se
rect 7616 8704 8024 8840
tri 8024 8704 8160 8840 sw
rect 7480 8296 8160 8704
tri 7480 8160 7616 8296 ne
rect 7616 8160 8024 8296
tri 8024 8160 8160 8296 nw
tri 8840 8704 8976 8840 se
rect 8976 8704 9384 8840
tri 9384 8704 9520 8840 sw
tri 9520 8704 9656 8840 se
rect 9656 8704 10064 8840
tri 10064 8704 10200 8840 sw
rect 8840 8296 10200 8704
tri 8840 8160 8976 8296 ne
tri 6664 8024 6800 8160 sw
tri 6800 8024 6936 8160 se
rect 6936 8024 7344 8160
tri 7344 8024 7480 8160 sw
rect 4760 7616 7480 8024
tri 4760 7480 4896 7616 ne
tri 2584 7344 2720 7480 sw
tri 2720 7344 2856 7480 se
rect 2856 7344 3264 7480
tri 3264 7344 3400 7480 sw
tri 3400 7344 3536 7480 se
rect 3536 7344 3944 7480
tri 3944 7344 4080 7480 sw
tri 4080 7344 4216 7480 se
rect 4216 7344 4624 7480
tri 4624 7344 4760 7480 sw
tri 4760 7344 4896 7480 se
rect 4896 7344 5304 7616
tri 5304 7480 5440 7616 nw
tri 5440 7480 5576 7616 ne
rect 5576 7480 5984 7616
tri 5984 7480 6120 7616 nw
tri 6120 7480 6256 7616 ne
tri 5304 7344 5440 7480 sw
rect 0 6936 5440 7344
tri 0 6800 136 6936 ne
rect 136 6800 544 6936
tri 544 6800 680 6936 nw
tri 680 6800 816 6936 ne
tri 680 6664 816 6800 se
rect 816 6664 1224 6936
tri 1224 6800 1360 6936 nw
tri 1360 6800 1496 6936 ne
tri 1224 6664 1360 6800 sw
tri 1360 6664 1496 6800 se
rect 1496 6664 1904 6936
tri 1904 6800 2040 6936 nw
tri 2040 6800 2176 6936 ne
rect 2176 6800 2584 6936
tri 2584 6800 2720 6936 nw
tri 2720 6800 2856 6936 ne
tri 1904 6664 2040 6800 sw
rect 680 6256 2040 6664
tri 680 6120 816 6256 ne
rect 816 6120 1224 6256
tri 1224 6120 1360 6256 nw
tri 1360 6120 1496 6256 ne
rect 1496 6120 1904 6256
tri 1904 6120 2040 6256 nw
tri 2720 6664 2856 6800 se
rect 2856 6664 3264 6936
tri 3264 6800 3400 6936 nw
tri 3400 6800 3536 6936 ne
rect 3536 6800 3944 6936
tri 3944 6800 4080 6936 nw
tri 4080 6800 4216 6936 ne
rect 4216 6800 4624 6936
tri 4624 6800 4760 6936 nw
tri 4760 6800 4896 6936 ne
tri 3264 6664 3400 6800 sw
rect 2720 6256 3400 6664
tri 2720 6120 2856 6256 ne
tri 0 5984 136 6120 se
rect 136 5984 544 6120
tri 544 5984 680 6120 sw
rect 0 5576 680 5984
tri 0 5440 136 5576 ne
rect 136 5440 544 5576
tri 544 5440 680 5576 nw
tri 2720 5984 2856 6120 se
rect 2856 5984 3264 6256
tri 3264 6120 3400 6256 nw
tri 4760 6664 4896 6800 se
rect 4896 6664 5304 6936
tri 5304 6800 5440 6936 nw
tri 6120 7344 6256 7480 se
rect 6256 7344 6664 7616
tri 6664 7480 6800 7616 nw
tri 6800 7480 6936 7616 ne
rect 6936 7480 7344 7616
tri 7344 7480 7480 7616 nw
tri 8840 8024 8976 8160 se
rect 8976 8024 9384 8296
tri 9384 8160 9520 8296 nw
tri 9520 8160 9656 8296 ne
rect 9656 8160 10064 8296
tri 10064 8160 10200 8296 nw
tri 10880 8704 11016 8840 se
rect 11016 8704 11424 8840
tri 11424 8704 11560 8840 sw
rect 10880 8296 11560 8704
tri 10880 8160 11016 8296 ne
rect 11016 8160 11424 8296
tri 11424 8160 11560 8296 nw
tri 9384 8024 9520 8160 sw
rect 8840 7616 9520 8024
tri 8840 7480 8976 7616 ne
tri 6664 7344 6800 7480 sw
rect 6120 6936 6800 7344
tri 6120 6800 6256 6936 ne
tri 5304 6664 5440 6800 sw
tri 5440 6664 5576 6800 se
rect 5576 6664 5984 6800
tri 5984 6664 6120 6800 sw
tri 6120 6664 6256 6800 se
rect 6256 6664 6664 6936
tri 6664 6800 6800 6936 nw
tri 6664 6664 6800 6800 sw
rect 4760 6256 6800 6664
tri 4760 6120 4896 6256 ne
rect 4896 6120 5304 6256
tri 5304 6120 5440 6256 nw
tri 5440 6120 5576 6256 ne
tri 3264 5984 3400 6120 sw
tri 3400 5984 3536 6120 se
rect 3536 5984 3944 6120
tri 3944 5984 4080 6120 sw
tri 4080 5984 4216 6120 se
rect 4216 5984 4624 6120
tri 4624 5984 4760 6120 sw
rect 2720 5576 4760 5984
tri 2720 5440 2856 5576 ne
rect 2856 5440 3264 5576
tri 3264 5440 3400 5576 nw
tri 3400 5440 3536 5576 ne
rect 3536 5440 3944 5576
tri 3944 5440 4080 5576 nw
tri 4080 5440 4216 5576 ne
rect 4216 5440 4624 5576
tri 4624 5440 4760 5576 nw
tri 5440 5984 5576 6120 se
rect 5576 5984 5984 6256
tri 5984 6120 6120 6256 nw
tri 6120 6120 6256 6256 ne
tri 5984 5984 6120 6120 sw
tri 6120 5984 6256 6120 se
rect 6256 5984 6664 6256
tri 6664 6120 6800 6256 nw
tri 6664 5984 6800 6120 sw
rect 5440 5576 6800 5984
tri 5440 5440 5576 5576 ne
tri 5440 5304 5576 5440 se
rect 5576 5304 5984 5576
tri 5984 5440 6120 5576 nw
tri 6120 5440 6256 5576 ne
rect 6256 5440 6664 5576
tri 6664 5440 6800 5576 nw
tri 7480 7344 7616 7480 se
rect 7616 7344 8024 7480
tri 8024 7344 8160 7480 sw
rect 7480 6936 8160 7344
tri 7480 6800 7616 6936 ne
tri 7480 6664 7616 6800 se
rect 7616 6664 8024 6936
tri 8024 6800 8160 6936 nw
tri 8840 7344 8976 7480 se
rect 8976 7344 9384 7616
tri 9384 7480 9520 7616 nw
tri 9384 7344 9520 7480 sw
rect 8840 6936 9520 7344
tri 8840 6800 8976 6936 ne
tri 8024 6664 8160 6800 sw
tri 8160 6664 8296 6800 se
rect 8296 6664 8704 6800
tri 8704 6664 8840 6800 sw
tri 8840 6664 8976 6800 se
rect 8976 6664 9384 6936
tri 9384 6800 9520 6936 nw
tri 10200 8024 10336 8160 se
rect 10336 8024 10744 8160
tri 10744 8024 10880 8160 sw
rect 10200 7616 10880 8024
tri 10200 7480 10336 7616 ne
tri 10200 7344 10336 7480 se
rect 10336 7344 10744 7616
tri 10744 7480 10880 7616 nw
tri 12240 8024 12376 8160 se
rect 12376 8024 12784 8160
tri 12784 8024 12920 8160 sw
rect 12240 7616 12920 8024
tri 12240 7480 12376 7616 ne
rect 12376 7480 12784 7616
tri 12784 7480 12920 7616 nw
tri 10744 7344 10880 7480 sw
tri 10880 7344 11016 7480 se
rect 11016 7344 11424 7480
tri 11424 7344 11560 7480 sw
tri 11560 7344 11696 7480 se
rect 11696 7344 12104 7480
tri 12104 7344 12240 7480 sw
rect 10200 6936 12240 7344
tri 10200 6800 10336 6936 ne
rect 10336 6800 10744 6936
tri 10744 6800 10880 6936 nw
tri 10880 6800 11016 6936 ne
rect 11016 6800 11424 6936
tri 11424 6800 11560 6936 nw
tri 11560 6800 11696 6936 ne
rect 11696 6800 12104 6936
tri 12104 6800 12240 6936 nw
tri 13600 7344 13736 7480 se
rect 13736 7344 14144 7480
tri 14144 7344 14280 7480 sw
rect 13600 6936 14280 7344
tri 13600 6800 13736 6936 ne
rect 13736 6800 14144 6936
tri 14144 6800 14280 6936 nw
tri 9384 6664 9520 6800 sw
tri 9520 6664 9656 6800 se
rect 9656 6664 10064 6800
tri 10064 6664 10200 6800 sw
rect 7480 6256 10200 6664
tri 7480 6120 7616 6256 ne
tri 7480 5984 7616 6120 se
rect 7616 5984 8024 6256
tri 8024 6120 8160 6256 nw
tri 8160 6120 8296 6256 ne
tri 8024 5984 8160 6120 sw
tri 8160 5984 8296 6120 se
rect 8296 5984 8704 6256
tri 8704 6120 8840 6256 nw
tri 8840 6120 8976 6256 ne
rect 8976 6120 9384 6256
tri 9384 6120 9520 6256 nw
tri 9520 6120 9656 6256 ne
rect 9656 6120 10064 6256
tri 10064 6120 10200 6256 nw
tri 12920 6664 13056 6800 se
rect 13056 6664 13464 6800
tri 13464 6664 13600 6800 sw
rect 12920 6256 13600 6664
tri 12920 6120 13056 6256 ne
rect 13056 6120 13464 6256
tri 13464 6120 13600 6256 nw
tri 8704 5984 8840 6120 sw
rect 7480 5576 8840 5984
tri 7480 5440 7616 5576 ne
tri 5984 5304 6120 5440 sw
rect 5440 4896 6120 5304
tri 5440 4760 5576 4896 ne
tri 0 4624 136 4760 se
rect 136 4624 544 4760
tri 544 4624 680 4760 sw
tri 680 4624 816 4760 se
rect 816 4624 1224 4760
tri 1224 4624 1360 4760 sw
tri 1360 4624 1496 4760 se
rect 1496 4624 1904 4760
tri 1904 4624 2040 4760 sw
tri 2040 4624 2176 4760 se
rect 2176 4624 2584 4760
tri 2584 4624 2720 4760 sw
tri 2720 4624 2856 4760 se
rect 2856 4624 3264 4760
tri 3264 4624 3400 4760 sw
tri 3400 4624 3536 4760 se
rect 3536 4624 3944 4760
tri 3944 4624 4080 4760 sw
tri 4080 4624 4216 4760 se
rect 4216 4624 4624 4760
tri 4624 4624 4760 4760 sw
rect 0 4216 4760 4624
tri 0 4080 136 4216 ne
tri 0 3944 136 4080 se
rect 136 3944 544 4216
tri 544 4080 680 4216 nw
tri 680 4080 816 4216 ne
rect 816 4080 1224 4216
tri 1224 4080 1360 4216 nw
tri 1360 4080 1496 4216 ne
rect 1496 4080 1904 4216
tri 1904 4080 2040 4216 nw
tri 2040 4080 2176 4216 ne
rect 2176 4080 2584 4216
tri 2584 4080 2720 4216 nw
tri 2720 4080 2856 4216 ne
rect 2856 4080 3264 4216
tri 3264 4080 3400 4216 nw
tri 3400 4080 3536 4216 ne
rect 3536 4080 3944 4216
tri 3944 4080 4080 4216 nw
tri 4080 4080 4216 4216 ne
tri 544 3944 680 4080 sw
rect 0 3536 680 3944
tri 0 3400 136 3536 ne
tri 0 3264 136 3400 se
rect 136 3264 544 3536
tri 544 3400 680 3536 nw
tri 4080 3944 4216 4080 se
rect 4216 3944 4624 4216
tri 4624 4080 4760 4216 nw
tri 5440 4624 5576 4760 se
rect 5576 4624 5984 4896
tri 5984 4760 6120 4896 nw
tri 6800 5304 6936 5440 se
rect 6936 5304 7344 5440
tri 7344 5304 7480 5440 sw
tri 7480 5304 7616 5440 se
rect 7616 5304 8024 5576
tri 8024 5440 8160 5576 nw
tri 8160 5440 8296 5576 ne
tri 8024 5304 8160 5440 sw
tri 8160 5304 8296 5440 se
rect 8296 5304 8704 5576
tri 8704 5440 8840 5576 nw
tri 10880 5984 11016 6120 se
rect 11016 5984 11424 6120
tri 11424 5984 11560 6120 sw
rect 10880 5576 11560 5984
tri 10880 5440 11016 5576 ne
rect 11016 5440 11424 5576
tri 11424 5440 11560 5576 nw
tri 12240 5984 12376 6120 se
rect 12376 5984 12784 6120
tri 12784 5984 12920 6120 sw
rect 12240 5576 12920 5984
tri 12240 5440 12376 5576 ne
rect 12376 5440 12784 5576
tri 12784 5440 12920 5576 nw
tri 8704 5304 8840 5440 sw
tri 8840 5304 8976 5440 se
rect 8976 5304 9384 5440
tri 9384 5304 9520 5440 sw
rect 6800 4896 9520 5304
tri 6800 4760 6936 4896 ne
tri 5984 4624 6120 4760 sw
tri 6120 4624 6256 4760 se
rect 6256 4624 6664 4760
tri 6664 4624 6800 4760 sw
tri 6800 4624 6936 4760 se
rect 6936 4624 7344 4896
tri 7344 4760 7480 4896 nw
tri 7480 4760 7616 4896 ne
tri 7344 4624 7480 4760 sw
tri 7480 4624 7616 4760 se
rect 7616 4624 8024 4896
tri 8024 4760 8160 4896 nw
tri 8160 4760 8296 4896 ne
tri 8024 4624 8160 4760 sw
tri 8160 4624 8296 4760 se
rect 8296 4624 8704 4896
tri 8704 4760 8840 4896 nw
tri 8840 4760 8976 4896 ne
rect 8976 4760 9384 4896
tri 9384 4760 9520 4896 nw
tri 10200 5304 10336 5440 se
rect 10336 5304 10744 5440
tri 10744 5304 10880 5440 sw
rect 10200 4896 10880 5304
tri 10200 4760 10336 4896 ne
rect 10336 4760 10744 4896
tri 10744 4760 10880 4896 nw
tri 11560 5304 11696 5440 se
rect 11696 5304 12104 5440
tri 12104 5304 12240 5440 sw
rect 11560 4896 12240 5304
tri 11560 4760 11696 4896 ne
rect 11696 4760 12104 4896
tri 12104 4760 12240 4896 nw
tri 13600 5304 13736 5440 se
rect 13736 5304 14144 5440
tri 14144 5304 14280 5440 sw
rect 13600 4896 14280 5304
tri 13600 4760 13736 4896 ne
rect 13736 4760 14144 4896
tri 14144 4760 14280 4896 nw
tri 8704 4624 8840 4760 sw
rect 5440 4216 8840 4624
tri 5440 4080 5576 4216 ne
rect 5576 4080 5984 4216
tri 5984 4080 6120 4216 nw
tri 6120 4080 6256 4216 ne
rect 6256 4080 6664 4216
tri 6664 4080 6800 4216 nw
tri 6800 4080 6936 4216 ne
rect 6936 4080 7344 4216
tri 7344 4080 7480 4216 nw
tri 7480 4080 7616 4216 ne
rect 7616 4080 8024 4216
tri 8024 4080 8160 4216 nw
tri 8160 4080 8296 4216 ne
rect 8296 4080 8704 4216
tri 8704 4080 8840 4216 nw
tri 10880 4624 11016 4760 se
rect 11016 4624 11424 4760
tri 11424 4624 11560 4760 sw
rect 10880 4216 11560 4624
tri 10880 4080 11016 4216 ne
rect 11016 4080 11424 4216
tri 11424 4080 11560 4216 nw
tri 12920 4624 13056 4760 se
rect 13056 4624 13464 4760
tri 13464 4624 13600 4760 sw
rect 12920 4216 13600 4624
tri 12920 4080 13056 4216 ne
rect 13056 4080 13464 4216
tri 13464 4080 13600 4216 nw
tri 4624 3944 4760 4080 sw
rect 4080 3536 4760 3944
tri 4080 3400 4216 3536 ne
tri 544 3264 680 3400 sw
rect 0 2856 680 3264
tri 0 2720 136 2856 ne
tri 0 2584 136 2720 se
rect 136 2584 544 2856
tri 544 2720 680 2856 nw
tri 544 2584 680 2720 sw
rect 0 2176 680 2584
tri 0 2040 136 2176 ne
tri 0 1904 136 2040 se
rect 136 1904 544 2176
tri 544 2040 680 2176 nw
tri 544 1904 680 2040 sw
rect 0 1496 680 1904
tri 0 1360 136 1496 ne
tri 0 1224 136 1360 se
rect 136 1224 544 1496
tri 544 1360 680 1496 nw
tri 1360 3264 1496 3400 se
rect 1496 3264 1904 3400
tri 1904 3264 2040 3400 sw
tri 2040 3264 2176 3400 se
rect 2176 3264 2584 3400
tri 2584 3264 2720 3400 sw
tri 2720 3264 2856 3400 se
rect 2856 3264 3264 3400
tri 3264 3264 3400 3400 sw
rect 1360 2856 3400 3264
tri 1360 2720 1496 2856 ne
tri 1360 2584 1496 2720 se
rect 1496 2584 1904 2856
tri 1904 2720 2040 2856 nw
tri 2040 2720 2176 2856 ne
tri 1904 2584 2040 2720 sw
tri 2040 2584 2176 2720 se
rect 2176 2584 2584 2856
tri 2584 2720 2720 2856 nw
tri 2720 2720 2856 2856 ne
tri 2584 2584 2720 2720 sw
tri 2720 2584 2856 2720 se
rect 2856 2584 3264 2856
tri 3264 2720 3400 2856 nw
tri 3264 2584 3400 2720 sw
rect 1360 2176 3400 2584
tri 1360 2040 1496 2176 ne
tri 1360 1904 1496 2040 se
rect 1496 1904 1904 2176
tri 1904 2040 2040 2176 nw
tri 2040 2040 2176 2176 ne
tri 1904 1904 2040 2040 sw
tri 2040 1904 2176 2040 se
rect 2176 1904 2584 2176
tri 2584 2040 2720 2176 nw
tri 2720 2040 2856 2176 ne
tri 2584 1904 2720 2040 sw
tri 2720 1904 2856 2040 se
rect 2856 1904 3264 2176
tri 3264 2040 3400 2176 nw
tri 3264 1904 3400 2040 sw
rect 1360 1496 3400 1904
tri 1360 1360 1496 1496 ne
rect 1496 1360 1904 1496
tri 1904 1360 2040 1496 nw
tri 2040 1360 2176 1496 ne
rect 2176 1360 2584 1496
tri 2584 1360 2720 1496 nw
tri 2720 1360 2856 1496 ne
rect 2856 1360 3264 1496
tri 3264 1360 3400 1496 nw
tri 4080 3264 4216 3400 se
rect 4216 3264 4624 3536
tri 4624 3400 4760 3536 nw
tri 9520 3944 9656 4080 se
rect 9656 3944 10064 4080
tri 10064 3944 10200 4080 sw
rect 9520 3536 10200 3944
tri 9520 3400 9656 3536 ne
tri 4624 3264 4760 3400 sw
rect 4080 2856 4760 3264
tri 4080 2720 4216 2856 ne
tri 4080 2584 4216 2720 se
rect 4216 2584 4624 2856
tri 4624 2720 4760 2856 nw
tri 6120 3264 6256 3400 se
rect 6256 3264 6664 3400
tri 6664 3264 6800 3400 sw
tri 6800 3264 6936 3400 se
rect 6936 3264 7344 3400
tri 7344 3264 7480 3400 sw
tri 7480 3264 7616 3400 se
rect 7616 3264 8024 3400
tri 8024 3264 8160 3400 sw
rect 6120 2856 8160 3264
tri 6120 2720 6256 2856 ne
rect 6256 2720 6664 2856
tri 6664 2720 6800 2856 nw
tri 6800 2720 6936 2856 ne
tri 4624 2584 4760 2720 sw
rect 4080 2176 4760 2584
tri 4080 2040 4216 2176 ne
tri 4080 1904 4216 2040 se
rect 4216 1904 4624 2176
tri 4624 2040 4760 2176 nw
tri 4624 1904 4760 2040 sw
rect 4080 1496 4760 1904
tri 4080 1360 4216 1496 ne
tri 544 1224 680 1360 sw
rect 0 816 680 1224
tri 0 680 136 816 ne
tri 0 544 136 680 se
rect 136 544 544 816
tri 544 680 680 816 nw
tri 4080 1224 4216 1360 se
rect 4216 1224 4624 1496
tri 4624 1360 4760 1496 nw
tri 5440 2584 5576 2720 se
rect 5576 2584 5984 2720
tri 5984 2584 6120 2720 sw
rect 5440 2176 6120 2584
tri 5440 2040 5576 2176 ne
tri 5440 1904 5576 2040 se
rect 5576 1904 5984 2176
tri 5984 2040 6120 2176 nw
tri 6800 2584 6936 2720 se
rect 6936 2584 7344 2856
tri 7344 2720 7480 2856 nw
tri 7480 2720 7616 2856 ne
rect 7616 2720 8024 2856
tri 8024 2720 8160 2856 nw
tri 9520 3264 9656 3400 se
rect 9656 3264 10064 3536
tri 10064 3400 10200 3536 nw
tri 12240 3944 12376 4080 se
rect 12376 3944 12784 4080
tri 12784 3944 12920 4080 sw
rect 12240 3536 12920 3944
tri 12240 3400 12376 3536 ne
rect 12376 3400 12784 3536
tri 12784 3400 12920 3536 nw
tri 13600 3944 13736 4080 se
rect 13736 3944 14144 4080
tri 14144 3944 14280 4080 sw
rect 13600 3536 14280 3944
tri 13600 3400 13736 3536 ne
tri 10064 3264 10200 3400 sw
rect 9520 2856 10200 3264
tri 9520 2720 9656 2856 ne
tri 7344 2584 7480 2720 sw
rect 6800 2176 7480 2584
tri 6800 2040 6936 2176 ne
rect 6936 2040 7344 2176
tri 7344 2040 7480 2176 nw
tri 8160 2584 8296 2720 se
rect 8296 2584 8704 2720
tri 8704 2584 8840 2720 sw
rect 8160 2176 8840 2584
tri 8160 2040 8296 2176 ne
rect 8296 2040 8704 2176
tri 8704 2040 8840 2176 nw
tri 9520 2584 9656 2720 se
rect 9656 2584 10064 2856
tri 10064 2720 10200 2856 nw
tri 11560 3264 11696 3400 se
rect 11696 3264 12104 3400
tri 12104 3264 12240 3400 sw
rect 11560 2856 12240 3264
tri 11560 2720 11696 2856 ne
rect 11696 2720 12104 2856
tri 12104 2720 12240 2856 nw
tri 13600 3264 13736 3400 se
rect 13736 3264 14144 3536
tri 14144 3400 14280 3536 nw
tri 14144 3264 14280 3400 sw
rect 13600 2856 14280 3264
tri 13600 2720 13736 2856 ne
rect 13736 2720 14144 2856
tri 14144 2720 14280 2856 nw
tri 10064 2584 10200 2720 sw
rect 9520 2176 10200 2584
tri 9520 2040 9656 2176 ne
rect 9656 2040 10064 2176
tri 10064 2040 10200 2176 nw
tri 10880 2584 11016 2720 se
rect 11016 2584 11424 2720
tri 11424 2584 11560 2720 sw
rect 10880 2176 11560 2584
tri 10880 2040 11016 2176 ne
tri 5984 1904 6120 2040 sw
rect 5440 1496 6120 1904
tri 5440 1360 5576 1496 ne
rect 5576 1360 5984 1496
tri 5984 1360 6120 1496 nw
tri 7480 1904 7616 2040 se
rect 7616 1904 8024 2040
tri 8024 1904 8160 2040 sw
rect 7480 1496 8160 1904
tri 7480 1360 7616 1496 ne
tri 4624 1224 4760 1360 sw
rect 4080 816 4760 1224
tri 4080 680 4216 816 ne
tri 544 544 680 680 sw
tri 680 544 816 680 se
rect 816 544 1224 680
tri 1224 544 1360 680 sw
tri 1360 544 1496 680 se
rect 1496 544 1904 680
tri 1904 544 2040 680 sw
tri 2040 544 2176 680 se
rect 2176 544 2584 680
tri 2584 544 2720 680 sw
tri 2720 544 2856 680 se
rect 2856 544 3264 680
tri 3264 544 3400 680 sw
tri 3400 544 3536 680 se
rect 3536 544 3944 680
tri 3944 544 4080 680 sw
tri 4080 544 4216 680 se
rect 4216 544 4624 816
tri 4624 680 4760 816 nw
tri 6120 1224 6256 1360 se
rect 6256 1224 6664 1360
tri 6664 1224 6800 1360 sw
tri 6800 1224 6936 1360 se
rect 6936 1224 7344 1360
tri 7344 1224 7480 1360 sw
tri 7480 1224 7616 1360 se
rect 7616 1224 8024 1496
tri 8024 1360 8160 1496 nw
tri 10880 1904 11016 2040 se
rect 11016 1904 11424 2176
tri 11424 2040 11560 2176 nw
tri 12920 2584 13056 2720 se
rect 13056 2584 13464 2720
tri 13464 2584 13600 2720 sw
rect 12920 2176 13600 2584
tri 12920 2040 13056 2176 ne
rect 13056 2040 13464 2176
tri 13464 2040 13600 2176 nw
tri 11424 1904 11560 2040 sw
rect 10880 1496 11560 1904
tri 10880 1360 11016 1496 ne
tri 8024 1224 8160 1360 sw
rect 6120 816 8160 1224
tri 6120 680 6256 816 ne
rect 6256 680 6664 816
tri 6664 680 6800 816 nw
tri 6800 680 6936 816 ne
rect 6936 680 7344 816
tri 7344 680 7480 816 nw
tri 7480 680 7616 816 ne
rect 7616 680 8024 816
tri 8024 680 8160 816 nw
tri 8840 1224 8976 1360 se
rect 8976 1224 9384 1360
tri 9384 1224 9520 1360 sw
rect 8840 816 9520 1224
tri 8840 680 8976 816 ne
rect 8976 680 9384 816
tri 9384 680 9520 816 nw
tri 10880 1224 11016 1360 se
rect 11016 1224 11424 1496
tri 11424 1360 11560 1496 nw
tri 12240 1904 12376 2040 se
rect 12376 1904 12784 2040
tri 12784 1904 12920 2040 sw
rect 12240 1496 12920 1904
tri 12240 1360 12376 1496 ne
rect 12376 1360 12784 1496
tri 12784 1360 12920 1496 nw
tri 11424 1224 11560 1360 sw
tri 11560 1224 11696 1360 se
rect 11696 1224 12104 1360
tri 12104 1224 12240 1360 sw
rect 10880 816 12240 1224
tri 10880 680 11016 816 ne
rect 11016 680 11424 816
tri 11424 680 11560 816 nw
tri 11560 680 11696 816 ne
rect 11696 680 12104 816
tri 12104 680 12240 816 nw
tri 12920 1224 13056 1360 se
rect 13056 1224 13464 1360
tri 13464 1224 13600 1360 sw
tri 13600 1224 13736 1360 se
rect 13736 1224 14144 1360
tri 14144 1224 14280 1360 sw
rect 12920 816 14280 1224
tri 12920 680 13056 816 ne
tri 4624 544 4760 680 sw
rect 0 136 4760 544
tri 0 0 136 136 ne
rect 136 0 544 136
tri 544 0 680 136 nw
tri 680 0 816 136 ne
rect 816 0 1224 136
tri 1224 0 1360 136 nw
tri 1360 0 1496 136 ne
rect 1496 0 1904 136
tri 1904 0 2040 136 nw
tri 2040 0 2176 136 ne
rect 2176 0 2584 136
tri 2584 0 2720 136 nw
tri 2720 0 2856 136 ne
rect 2856 0 3264 136
tri 3264 0 3400 136 nw
tri 3400 0 3536 136 ne
rect 3536 0 3944 136
tri 3944 0 4080 136 nw
tri 4080 0 4216 136 ne
rect 4216 0 4624 136
tri 4624 0 4760 136 nw
tri 8160 544 8296 680 se
rect 8296 544 8704 680
tri 8704 544 8840 680 sw
rect 8160 136 8840 544
tri 8160 0 8296 136 ne
rect 8296 0 8704 136
tri 8704 0 8840 136 nw
tri 10200 544 10336 680 se
rect 10336 544 10744 680
tri 10744 544 10880 680 sw
rect 10200 136 10880 544
tri 10200 0 10336 136 ne
rect 10336 0 10744 136
tri 10744 0 10880 136 nw
tri 12920 544 13056 680 se
rect 13056 544 13464 816
tri 13464 680 13600 816 nw
tri 13600 680 13736 816 ne
rect 13736 680 14144 816
tri 14144 680 14280 816 nw
tri 13464 544 13600 680 sw
rect 12920 136 13600 544
tri 12920 0 13056 136 ne
rect 13056 0 13464 136
tri 13464 0 13600 136 nw
<< metal4 >>
tri 0 14144 136 14280 se
rect 136 14144 544 14280
tri 544 14144 680 14280 sw
tri 680 14144 816 14280 se
rect 816 14144 1224 14280
tri 1224 14144 1360 14280 sw
tri 1360 14144 1496 14280 se
rect 1496 14144 1904 14280
tri 1904 14144 2040 14280 sw
tri 2040 14144 2176 14280 se
rect 2176 14144 2584 14280
tri 2584 14144 2720 14280 sw
tri 2720 14144 2856 14280 se
rect 2856 14144 3264 14280
tri 3264 14144 3400 14280 sw
tri 3400 14144 3536 14280 se
rect 3536 14144 3944 14280
tri 3944 14144 4080 14280 sw
tri 4080 14144 4216 14280 se
rect 4216 14144 4624 14280
tri 4624 14144 4760 14280 sw
rect 0 13736 4760 14144
tri 0 13600 136 13736 ne
tri 0 13464 136 13600 se
rect 136 13464 544 13736
tri 544 13600 680 13736 nw
tri 680 13600 816 13736 ne
rect 816 13600 1224 13736
tri 1224 13600 1360 13736 nw
tri 1360 13600 1496 13736 ne
rect 1496 13600 1904 13736
tri 1904 13600 2040 13736 nw
tri 2040 13600 2176 13736 ne
rect 2176 13600 2584 13736
tri 2584 13600 2720 13736 nw
tri 2720 13600 2856 13736 ne
rect 2856 13600 3264 13736
tri 3264 13600 3400 13736 nw
tri 3400 13600 3536 13736 ne
rect 3536 13600 3944 13736
tri 3944 13600 4080 13736 nw
tri 4080 13600 4216 13736 ne
tri 544 13464 680 13600 sw
rect 0 13056 680 13464
tri 0 12920 136 13056 ne
tri 0 12784 136 12920 se
rect 136 12784 544 13056
tri 544 12920 680 13056 nw
tri 4080 13464 4216 13600 se
rect 4216 13464 4624 13736
tri 4624 13600 4760 13736 nw
tri 6120 14144 6256 14280 se
rect 6256 14144 6664 14280
tri 6664 14144 6800 14280 sw
tri 6800 14144 6936 14280 se
rect 6936 14144 7344 14280
tri 7344 14144 7480 14280 sw
rect 6120 13736 7480 14144
tri 6120 13600 6256 13736 ne
rect 6256 13600 6664 13736
tri 6664 13600 6800 13736 nw
tri 6800 13600 6936 13736 ne
tri 4624 13464 4760 13600 sw
rect 4080 13056 4760 13464
tri 4080 12920 4216 13056 ne
tri 544 12784 680 12920 sw
rect 0 12376 680 12784
tri 0 12240 136 12376 ne
tri 0 12104 136 12240 se
rect 136 12104 544 12376
tri 544 12240 680 12376 nw
tri 544 12104 680 12240 sw
rect 0 11696 680 12104
tri 0 11560 136 11696 ne
tri 0 11424 136 11560 se
rect 136 11424 544 11696
tri 544 11560 680 11696 nw
tri 544 11424 680 11560 sw
rect 0 11016 680 11424
tri 0 10880 136 11016 ne
tri 0 10744 136 10880 se
rect 136 10744 544 11016
tri 544 10880 680 11016 nw
tri 1360 12784 1496 12920 se
rect 1496 12784 1904 12920
tri 1904 12784 2040 12920 sw
tri 2040 12784 2176 12920 se
rect 2176 12784 2584 12920
tri 2584 12784 2720 12920 sw
tri 2720 12784 2856 12920 se
rect 2856 12784 3264 12920
tri 3264 12784 3400 12920 sw
rect 1360 12376 3400 12784
tri 1360 12240 1496 12376 ne
tri 1360 12104 1496 12240 se
rect 1496 12104 1904 12376
tri 1904 12240 2040 12376 nw
tri 2040 12240 2176 12376 ne
tri 1904 12104 2040 12240 sw
tri 2040 12104 2176 12240 se
rect 2176 12104 2584 12376
tri 2584 12240 2720 12376 nw
tri 2720 12240 2856 12376 ne
tri 2584 12104 2720 12240 sw
tri 2720 12104 2856 12240 se
rect 2856 12104 3264 12376
tri 3264 12240 3400 12376 nw
tri 3264 12104 3400 12240 sw
rect 1360 11696 3400 12104
tri 1360 11560 1496 11696 ne
tri 1360 11424 1496 11560 se
rect 1496 11424 1904 11696
tri 1904 11560 2040 11696 nw
tri 2040 11560 2176 11696 ne
tri 1904 11424 2040 11560 sw
tri 2040 11424 2176 11560 se
rect 2176 11424 2584 11696
tri 2584 11560 2720 11696 nw
tri 2720 11560 2856 11696 ne
tri 2584 11424 2720 11560 sw
tri 2720 11424 2856 11560 se
rect 2856 11424 3264 11696
tri 3264 11560 3400 11696 nw
tri 3264 11424 3400 11560 sw
rect 1360 11016 3400 11424
tri 1360 10880 1496 11016 ne
rect 1496 10880 1904 11016
tri 1904 10880 2040 11016 nw
tri 2040 10880 2176 11016 ne
rect 2176 10880 2584 11016
tri 2584 10880 2720 11016 nw
tri 2720 10880 2856 11016 ne
rect 2856 10880 3264 11016
tri 3264 10880 3400 11016 nw
tri 4080 12784 4216 12920 se
rect 4216 12784 4624 13056
tri 4624 12920 4760 13056 nw
tri 6800 13464 6936 13600 se
rect 6936 13464 7344 13736
tri 7344 13600 7480 13736 nw
tri 8160 14144 8296 14280 se
rect 8296 14144 8704 14280
tri 8704 14144 8840 14280 sw
rect 8160 13736 8840 14144
tri 8160 13600 8296 13736 ne
rect 8296 13600 8704 13736
tri 8704 13600 8840 13736 nw
tri 9520 14144 9656 14280 se
rect 9656 14144 10064 14280
tri 10064 14144 10200 14280 sw
tri 10200 14144 10336 14280 se
rect 10336 14144 10744 14280
tri 10744 14144 10880 14280 sw
tri 10880 14144 11016 14280 se
rect 11016 14144 11424 14280
tri 11424 14144 11560 14280 sw
tri 11560 14144 11696 14280 se
rect 11696 14144 12104 14280
tri 12104 14144 12240 14280 sw
tri 12240 14144 12376 14280 se
rect 12376 14144 12784 14280
tri 12784 14144 12920 14280 sw
tri 12920 14144 13056 14280 se
rect 13056 14144 13464 14280
tri 13464 14144 13600 14280 sw
tri 13600 14144 13736 14280 se
rect 13736 14144 14144 14280
tri 14144 14144 14280 14280 sw
rect 9520 13736 14280 14144
tri 9520 13600 9656 13736 ne
tri 7344 13464 7480 13600 sw
tri 7480 13464 7616 13600 se
rect 7616 13464 8024 13600
tri 8024 13464 8160 13600 sw
rect 6800 13056 8160 13464
tri 6800 12920 6936 13056 ne
rect 6936 12920 7344 13056
tri 7344 12920 7480 13056 nw
tri 7480 12920 7616 13056 ne
tri 4624 12784 4760 12920 sw
rect 4080 12376 4760 12784
tri 4080 12240 4216 12376 ne
tri 4080 12104 4216 12240 se
rect 4216 12104 4624 12376
tri 4624 12240 4760 12376 nw
tri 7480 12784 7616 12920 se
rect 7616 12784 8024 13056
tri 8024 12920 8160 13056 nw
tri 9520 13464 9656 13600 se
rect 9656 13464 10064 13736
tri 10064 13600 10200 13736 nw
tri 10200 13600 10336 13736 ne
rect 10336 13600 10744 13736
tri 10744 13600 10880 13736 nw
tri 10880 13600 11016 13736 ne
rect 11016 13600 11424 13736
tri 11424 13600 11560 13736 nw
tri 11560 13600 11696 13736 ne
rect 11696 13600 12104 13736
tri 12104 13600 12240 13736 nw
tri 12240 13600 12376 13736 ne
rect 12376 13600 12784 13736
tri 12784 13600 12920 13736 nw
tri 12920 13600 13056 13736 ne
rect 13056 13600 13464 13736
tri 13464 13600 13600 13736 nw
tri 13600 13600 13736 13736 ne
tri 10064 13464 10200 13600 sw
rect 9520 13056 10200 13464
tri 9520 12920 9656 13056 ne
tri 8024 12784 8160 12920 sw
tri 8160 12784 8296 12920 se
rect 8296 12784 8704 12920
tri 8704 12784 8840 12920 sw
rect 7480 12376 8840 12784
tri 7480 12240 7616 12376 ne
tri 4624 12104 4760 12240 sw
rect 4080 11696 4760 12104
tri 4080 11560 4216 11696 ne
tri 4080 11424 4216 11560 se
rect 4216 11424 4624 11696
tri 4624 11560 4760 11696 nw
tri 6120 12104 6256 12240 se
rect 6256 12104 6664 12240
tri 6664 12104 6800 12240 sw
rect 6120 11696 6800 12104
tri 6120 11560 6256 11696 ne
tri 4624 11424 4760 11560 sw
rect 4080 11016 4760 11424
tri 4080 10880 4216 11016 ne
tri 544 10744 680 10880 sw
rect 0 10336 680 10744
tri 0 10200 136 10336 ne
tri 0 10064 136 10200 se
rect 136 10064 544 10336
tri 544 10200 680 10336 nw
tri 4080 10744 4216 10880 se
rect 4216 10744 4624 11016
tri 4624 10880 4760 11016 nw
tri 5440 11424 5576 11560 se
rect 5576 11424 5984 11560
tri 5984 11424 6120 11560 sw
tri 6120 11424 6256 11560 se
rect 6256 11424 6664 11696
tri 6664 11560 6800 11696 nw
tri 7480 12104 7616 12240 se
rect 7616 12104 8024 12376
tri 8024 12240 8160 12376 nw
tri 8160 12240 8296 12376 ne
tri 8024 12104 8160 12240 sw
tri 8160 12104 8296 12240 se
rect 8296 12104 8704 12376
tri 8704 12240 8840 12376 nw
tri 8704 12104 8840 12240 sw
rect 7480 11696 8840 12104
tri 7480 11560 7616 11696 ne
rect 7616 11560 8024 11696
tri 8024 11560 8160 11696 nw
tri 8160 11560 8296 11696 ne
rect 8296 11560 8704 11696
tri 8704 11560 8840 11696 nw
tri 9520 12784 9656 12920 se
rect 9656 12784 10064 13056
tri 10064 12920 10200 13056 nw
tri 13600 13464 13736 13600 se
rect 13736 13464 14144 13736
tri 14144 13600 14280 13736 nw
tri 14144 13464 14280 13600 sw
rect 13600 13056 14280 13464
tri 13600 12920 13736 13056 ne
tri 10064 12784 10200 12920 sw
rect 9520 12376 10200 12784
tri 9520 12240 9656 12376 ne
tri 9520 12104 9656 12240 se
rect 9656 12104 10064 12376
tri 10064 12240 10200 12376 nw
tri 10064 12104 10200 12240 sw
rect 9520 11696 10200 12104
tri 9520 11560 9656 11696 ne
tri 6664 11424 6800 11560 sw
rect 5440 11016 6800 11424
tri 5440 10880 5576 11016 ne
rect 5576 10880 5984 11016
tri 5984 10880 6120 11016 nw
tri 6120 10880 6256 11016 ne
tri 4624 10744 4760 10880 sw
rect 4080 10336 4760 10744
tri 4080 10200 4216 10336 ne
tri 544 10064 680 10200 sw
tri 680 10064 816 10200 se
rect 816 10064 1224 10200
tri 1224 10064 1360 10200 sw
tri 1360 10064 1496 10200 se
rect 1496 10064 1904 10200
tri 1904 10064 2040 10200 sw
tri 2040 10064 2176 10200 se
rect 2176 10064 2584 10200
tri 2584 10064 2720 10200 sw
tri 2720 10064 2856 10200 se
rect 2856 10064 3264 10200
tri 3264 10064 3400 10200 sw
tri 3400 10064 3536 10200 se
rect 3536 10064 3944 10200
tri 3944 10064 4080 10200 sw
tri 4080 10064 4216 10200 se
rect 4216 10064 4624 10336
tri 4624 10200 4760 10336 nw
tri 6120 10744 6256 10880 se
rect 6256 10744 6664 11016
tri 6664 10880 6800 11016 nw
tri 9520 11424 9656 11560 se
rect 9656 11424 10064 11696
tri 10064 11560 10200 11696 nw
tri 10064 11424 10200 11560 sw
rect 9520 11016 10200 11424
tri 9520 10880 9656 11016 ne
tri 6664 10744 6800 10880 sw
tri 6800 10744 6936 10880 se
rect 6936 10744 7344 10880
tri 7344 10744 7480 10880 sw
rect 6120 10336 7480 10744
tri 6120 10200 6256 10336 ne
rect 6256 10200 6664 10336
tri 6664 10200 6800 10336 nw
tri 6800 10200 6936 10336 ne
tri 4624 10064 4760 10200 sw
rect 0 9656 4760 10064
tri 0 9520 136 9656 ne
rect 136 9520 544 9656
tri 544 9520 680 9656 nw
tri 680 9520 816 9656 ne
rect 816 9520 1224 9656
tri 1224 9520 1360 9656 nw
tri 1360 9520 1496 9656 ne
rect 1496 9520 1904 9656
tri 1904 9520 2040 9656 nw
tri 2040 9520 2176 9656 ne
rect 2176 9520 2584 9656
tri 2584 9520 2720 9656 nw
tri 2720 9520 2856 9656 ne
rect 2856 9520 3264 9656
tri 3264 9520 3400 9656 nw
tri 3400 9520 3536 9656 ne
rect 3536 9520 3944 9656
tri 3944 9520 4080 9656 nw
tri 4080 9520 4216 9656 ne
rect 4216 9520 4624 9656
tri 4624 9520 4760 9656 nw
tri 5440 10064 5576 10200 se
rect 5576 10064 5984 10200
tri 5984 10064 6120 10200 sw
rect 5440 9656 6120 10064
tri 5440 9520 5576 9656 ne
tri 5440 9384 5576 9520 se
rect 5576 9384 5984 9656
tri 5984 9520 6120 9656 nw
tri 6800 10064 6936 10200 se
rect 6936 10064 7344 10336
tri 7344 10200 7480 10336 nw
tri 7344 10064 7480 10200 sw
rect 6800 9656 7480 10064
tri 6800 9520 6936 9656 ne
tri 5984 9384 6120 9520 sw
tri 6120 9384 6256 9520 se
rect 6256 9384 6664 9520
tri 6664 9384 6800 9520 sw
tri 6800 9384 6936 9520 se
rect 6936 9384 7344 9656
tri 7344 9520 7480 9656 nw
tri 8160 10744 8296 10880 se
rect 8296 10744 8704 10880
tri 8704 10744 8840 10880 sw
rect 8160 10336 8840 10744
tri 8160 10200 8296 10336 ne
tri 8160 10064 8296 10200 se
rect 8296 10064 8704 10336
tri 8704 10200 8840 10336 nw
tri 8704 10064 8840 10200 sw
rect 8160 9656 8840 10064
tri 8160 9520 8296 9656 ne
rect 8296 9520 8704 9656
tri 8704 9520 8840 9656 nw
tri 9520 10744 9656 10880 se
rect 9656 10744 10064 11016
tri 10064 10880 10200 11016 nw
tri 10880 12784 11016 12920 se
rect 11016 12784 11424 12920
tri 11424 12784 11560 12920 sw
tri 11560 12784 11696 12920 se
rect 11696 12784 12104 12920
tri 12104 12784 12240 12920 sw
tri 12240 12784 12376 12920 se
rect 12376 12784 12784 12920
tri 12784 12784 12920 12920 sw
rect 10880 12376 12920 12784
tri 10880 12240 11016 12376 ne
tri 10880 12104 11016 12240 se
rect 11016 12104 11424 12376
tri 11424 12240 11560 12376 nw
tri 11560 12240 11696 12376 ne
tri 11424 12104 11560 12240 sw
tri 11560 12104 11696 12240 se
rect 11696 12104 12104 12376
tri 12104 12240 12240 12376 nw
tri 12240 12240 12376 12376 ne
tri 12104 12104 12240 12240 sw
tri 12240 12104 12376 12240 se
rect 12376 12104 12784 12376
tri 12784 12240 12920 12376 nw
tri 12784 12104 12920 12240 sw
rect 10880 11696 12920 12104
tri 10880 11560 11016 11696 ne
tri 10880 11424 11016 11560 se
rect 11016 11424 11424 11696
tri 11424 11560 11560 11696 nw
tri 11560 11560 11696 11696 ne
tri 11424 11424 11560 11560 sw
tri 11560 11424 11696 11560 se
rect 11696 11424 12104 11696
tri 12104 11560 12240 11696 nw
tri 12240 11560 12376 11696 ne
tri 12104 11424 12240 11560 sw
tri 12240 11424 12376 11560 se
rect 12376 11424 12784 11696
tri 12784 11560 12920 11696 nw
tri 12784 11424 12920 11560 sw
rect 10880 11016 12920 11424
tri 10880 10880 11016 11016 ne
rect 11016 10880 11424 11016
tri 11424 10880 11560 11016 nw
tri 11560 10880 11696 11016 ne
rect 11696 10880 12104 11016
tri 12104 10880 12240 11016 nw
tri 12240 10880 12376 11016 ne
rect 12376 10880 12784 11016
tri 12784 10880 12920 11016 nw
tri 13600 12784 13736 12920 se
rect 13736 12784 14144 13056
tri 14144 12920 14280 13056 nw
tri 14144 12784 14280 12920 sw
rect 13600 12376 14280 12784
tri 13600 12240 13736 12376 ne
tri 13600 12104 13736 12240 se
rect 13736 12104 14144 12376
tri 14144 12240 14280 12376 nw
tri 14144 12104 14280 12240 sw
rect 13600 11696 14280 12104
tri 13600 11560 13736 11696 ne
tri 13600 11424 13736 11560 se
rect 13736 11424 14144 11696
tri 14144 11560 14280 11696 nw
tri 14144 11424 14280 11560 sw
rect 13600 11016 14280 11424
tri 13600 10880 13736 11016 ne
tri 10064 10744 10200 10880 sw
rect 9520 10336 10200 10744
tri 9520 10200 9656 10336 ne
tri 9520 10064 9656 10200 se
rect 9656 10064 10064 10336
tri 10064 10200 10200 10336 nw
tri 13600 10744 13736 10880 se
rect 13736 10744 14144 11016
tri 14144 10880 14280 11016 nw
tri 14144 10744 14280 10880 sw
rect 13600 10336 14280 10744
tri 13600 10200 13736 10336 ne
tri 10064 10064 10200 10200 sw
tri 10200 10064 10336 10200 se
rect 10336 10064 10744 10200
tri 10744 10064 10880 10200 sw
tri 10880 10064 11016 10200 se
rect 11016 10064 11424 10200
tri 11424 10064 11560 10200 sw
tri 11560 10064 11696 10200 se
rect 11696 10064 12104 10200
tri 12104 10064 12240 10200 sw
tri 12240 10064 12376 10200 se
rect 12376 10064 12784 10200
tri 12784 10064 12920 10200 sw
tri 12920 10064 13056 10200 se
rect 13056 10064 13464 10200
tri 13464 10064 13600 10200 sw
tri 13600 10064 13736 10200 se
rect 13736 10064 14144 10336
tri 14144 10200 14280 10336 nw
tri 14144 10064 14280 10200 sw
rect 9520 9656 14280 10064
tri 9520 9520 9656 9656 ne
rect 9656 9520 10064 9656
tri 10064 9520 10200 9656 nw
tri 10200 9520 10336 9656 ne
rect 10336 9520 10744 9656
tri 10744 9520 10880 9656 nw
tri 10880 9520 11016 9656 ne
rect 11016 9520 11424 9656
tri 11424 9520 11560 9656 nw
tri 11560 9520 11696 9656 ne
rect 11696 9520 12104 9656
tri 12104 9520 12240 9656 nw
tri 12240 9520 12376 9656 ne
rect 12376 9520 12784 9656
tri 12784 9520 12920 9656 nw
tri 12920 9520 13056 9656 ne
rect 13056 9520 13464 9656
tri 13464 9520 13600 9656 nw
tri 13600 9520 13736 9656 ne
rect 13736 9520 14144 9656
tri 14144 9520 14280 9656 nw
tri 7344 9384 7480 9520 sw
rect 5440 8976 7480 9384
tri 5440 8840 5576 8976 ne
tri 1360 8704 1496 8840 se
rect 1496 8704 1904 8840
tri 1904 8704 2040 8840 sw
tri 2040 8704 2176 8840 se
rect 2176 8704 2584 8840
tri 2584 8704 2720 8840 sw
rect 1360 8296 2720 8704
tri 1360 8160 1496 8296 ne
tri 1360 8024 1496 8160 se
rect 1496 8024 1904 8296
tri 1904 8160 2040 8296 nw
tri 2040 8160 2176 8296 ne
tri 1904 8024 2040 8160 sw
tri 2040 8024 2176 8160 se
rect 2176 8024 2584 8296
tri 2584 8160 2720 8296 nw
tri 4080 8704 4216 8840 se
rect 4216 8704 4624 8840
tri 4624 8704 4760 8840 sw
tri 4760 8704 4896 8840 se
rect 4896 8704 5304 8840
tri 5304 8704 5440 8840 sw
tri 5440 8704 5576 8840 se
rect 5576 8704 5984 8976
tri 5984 8840 6120 8976 nw
tri 6120 8840 6256 8976 ne
tri 5984 8704 6120 8840 sw
tri 6120 8704 6256 8840 se
rect 6256 8704 6664 8976
tri 6664 8840 6800 8976 nw
tri 6800 8840 6936 8976 ne
rect 6936 8840 7344 8976
tri 7344 8840 7480 8976 nw
tri 6664 8704 6800 8840 sw
rect 4080 8296 6800 8704
tri 4080 8160 4216 8296 ne
rect 4216 8160 4624 8296
tri 4624 8160 4760 8296 nw
tri 4760 8160 4896 8296 ne
tri 2584 8024 2720 8160 sw
rect 1360 7616 2720 8024
tri 1360 7480 1496 7616 ne
tri 0 7344 136 7480 se
rect 136 7344 544 7480
tri 544 7344 680 7480 sw
tri 680 7344 816 7480 se
rect 816 7344 1224 7480
tri 1224 7344 1360 7480 sw
tri 1360 7344 1496 7480 se
rect 1496 7344 1904 7616
tri 1904 7480 2040 7616 nw
tri 2040 7480 2176 7616 ne
tri 1904 7344 2040 7480 sw
tri 2040 7344 2176 7480 se
rect 2176 7344 2584 7616
tri 2584 7480 2720 7616 nw
tri 4760 8024 4896 8160 se
rect 4896 8024 5304 8296
tri 5304 8160 5440 8296 nw
tri 5440 8160 5576 8296 ne
tri 5304 8024 5440 8160 sw
tri 5440 8024 5576 8160 se
rect 5576 8024 5984 8296
tri 5984 8160 6120 8296 nw
tri 6120 8160 6256 8296 ne
tri 5984 8024 6120 8160 sw
tri 6120 8024 6256 8160 se
rect 6256 8024 6664 8296
tri 6664 8160 6800 8296 nw
tri 7480 8704 7616 8840 se
rect 7616 8704 8024 8840
tri 8024 8704 8160 8840 sw
rect 7480 8296 8160 8704
tri 7480 8160 7616 8296 ne
rect 7616 8160 8024 8296
tri 8024 8160 8160 8296 nw
tri 8840 8704 8976 8840 se
rect 8976 8704 9384 8840
tri 9384 8704 9520 8840 sw
tri 9520 8704 9656 8840 se
rect 9656 8704 10064 8840
tri 10064 8704 10200 8840 sw
rect 8840 8296 10200 8704
tri 8840 8160 8976 8296 ne
tri 6664 8024 6800 8160 sw
tri 6800 8024 6936 8160 se
rect 6936 8024 7344 8160
tri 7344 8024 7480 8160 sw
rect 4760 7616 7480 8024
tri 4760 7480 4896 7616 ne
tri 2584 7344 2720 7480 sw
tri 2720 7344 2856 7480 se
rect 2856 7344 3264 7480
tri 3264 7344 3400 7480 sw
tri 3400 7344 3536 7480 se
rect 3536 7344 3944 7480
tri 3944 7344 4080 7480 sw
tri 4080 7344 4216 7480 se
rect 4216 7344 4624 7480
tri 4624 7344 4760 7480 sw
tri 4760 7344 4896 7480 se
rect 4896 7344 5304 7616
tri 5304 7480 5440 7616 nw
tri 5440 7480 5576 7616 ne
rect 5576 7480 5984 7616
tri 5984 7480 6120 7616 nw
tri 6120 7480 6256 7616 ne
tri 5304 7344 5440 7480 sw
rect 0 6936 5440 7344
tri 0 6800 136 6936 ne
rect 136 6800 544 6936
tri 544 6800 680 6936 nw
tri 680 6800 816 6936 ne
tri 680 6664 816 6800 se
rect 816 6664 1224 6936
tri 1224 6800 1360 6936 nw
tri 1360 6800 1496 6936 ne
tri 1224 6664 1360 6800 sw
tri 1360 6664 1496 6800 se
rect 1496 6664 1904 6936
tri 1904 6800 2040 6936 nw
tri 2040 6800 2176 6936 ne
rect 2176 6800 2584 6936
tri 2584 6800 2720 6936 nw
tri 2720 6800 2856 6936 ne
tri 1904 6664 2040 6800 sw
rect 680 6256 2040 6664
tri 680 6120 816 6256 ne
rect 816 6120 1224 6256
tri 1224 6120 1360 6256 nw
tri 1360 6120 1496 6256 ne
rect 1496 6120 1904 6256
tri 1904 6120 2040 6256 nw
tri 2720 6664 2856 6800 se
rect 2856 6664 3264 6936
tri 3264 6800 3400 6936 nw
tri 3400 6800 3536 6936 ne
rect 3536 6800 3944 6936
tri 3944 6800 4080 6936 nw
tri 4080 6800 4216 6936 ne
rect 4216 6800 4624 6936
tri 4624 6800 4760 6936 nw
tri 4760 6800 4896 6936 ne
tri 3264 6664 3400 6800 sw
rect 2720 6256 3400 6664
tri 2720 6120 2856 6256 ne
tri 0 5984 136 6120 se
rect 136 5984 544 6120
tri 544 5984 680 6120 sw
rect 0 5576 680 5984
tri 0 5440 136 5576 ne
rect 136 5440 544 5576
tri 544 5440 680 5576 nw
tri 2720 5984 2856 6120 se
rect 2856 5984 3264 6256
tri 3264 6120 3400 6256 nw
tri 4760 6664 4896 6800 se
rect 4896 6664 5304 6936
tri 5304 6800 5440 6936 nw
tri 6120 7344 6256 7480 se
rect 6256 7344 6664 7616
tri 6664 7480 6800 7616 nw
tri 6800 7480 6936 7616 ne
rect 6936 7480 7344 7616
tri 7344 7480 7480 7616 nw
tri 8840 8024 8976 8160 se
rect 8976 8024 9384 8296
tri 9384 8160 9520 8296 nw
tri 9520 8160 9656 8296 ne
rect 9656 8160 10064 8296
tri 10064 8160 10200 8296 nw
tri 10880 8704 11016 8840 se
rect 11016 8704 11424 8840
tri 11424 8704 11560 8840 sw
rect 10880 8296 11560 8704
tri 10880 8160 11016 8296 ne
rect 11016 8160 11424 8296
tri 11424 8160 11560 8296 nw
tri 9384 8024 9520 8160 sw
rect 8840 7616 9520 8024
tri 8840 7480 8976 7616 ne
tri 6664 7344 6800 7480 sw
rect 6120 6936 6800 7344
tri 6120 6800 6256 6936 ne
tri 5304 6664 5440 6800 sw
tri 5440 6664 5576 6800 se
rect 5576 6664 5984 6800
tri 5984 6664 6120 6800 sw
tri 6120 6664 6256 6800 se
rect 6256 6664 6664 6936
tri 6664 6800 6800 6936 nw
tri 6664 6664 6800 6800 sw
rect 4760 6256 6800 6664
tri 4760 6120 4896 6256 ne
rect 4896 6120 5304 6256
tri 5304 6120 5440 6256 nw
tri 5440 6120 5576 6256 ne
tri 3264 5984 3400 6120 sw
tri 3400 5984 3536 6120 se
rect 3536 5984 3944 6120
tri 3944 5984 4080 6120 sw
tri 4080 5984 4216 6120 se
rect 4216 5984 4624 6120
tri 4624 5984 4760 6120 sw
rect 2720 5576 4760 5984
tri 2720 5440 2856 5576 ne
rect 2856 5440 3264 5576
tri 3264 5440 3400 5576 nw
tri 3400 5440 3536 5576 ne
rect 3536 5440 3944 5576
tri 3944 5440 4080 5576 nw
tri 4080 5440 4216 5576 ne
rect 4216 5440 4624 5576
tri 4624 5440 4760 5576 nw
tri 5440 5984 5576 6120 se
rect 5576 5984 5984 6256
tri 5984 6120 6120 6256 nw
tri 6120 6120 6256 6256 ne
tri 5984 5984 6120 6120 sw
tri 6120 5984 6256 6120 se
rect 6256 5984 6664 6256
tri 6664 6120 6800 6256 nw
tri 6664 5984 6800 6120 sw
rect 5440 5576 6800 5984
tri 5440 5440 5576 5576 ne
tri 5440 5304 5576 5440 se
rect 5576 5304 5984 5576
tri 5984 5440 6120 5576 nw
tri 6120 5440 6256 5576 ne
rect 6256 5440 6664 5576
tri 6664 5440 6800 5576 nw
tri 7480 7344 7616 7480 se
rect 7616 7344 8024 7480
tri 8024 7344 8160 7480 sw
rect 7480 6936 8160 7344
tri 7480 6800 7616 6936 ne
tri 7480 6664 7616 6800 se
rect 7616 6664 8024 6936
tri 8024 6800 8160 6936 nw
tri 8840 7344 8976 7480 se
rect 8976 7344 9384 7616
tri 9384 7480 9520 7616 nw
tri 9384 7344 9520 7480 sw
rect 8840 6936 9520 7344
tri 8840 6800 8976 6936 ne
tri 8024 6664 8160 6800 sw
tri 8160 6664 8296 6800 se
rect 8296 6664 8704 6800
tri 8704 6664 8840 6800 sw
tri 8840 6664 8976 6800 se
rect 8976 6664 9384 6936
tri 9384 6800 9520 6936 nw
tri 10200 8024 10336 8160 se
rect 10336 8024 10744 8160
tri 10744 8024 10880 8160 sw
rect 10200 7616 10880 8024
tri 10200 7480 10336 7616 ne
tri 10200 7344 10336 7480 se
rect 10336 7344 10744 7616
tri 10744 7480 10880 7616 nw
tri 12240 8024 12376 8160 se
rect 12376 8024 12784 8160
tri 12784 8024 12920 8160 sw
rect 12240 7616 12920 8024
tri 12240 7480 12376 7616 ne
rect 12376 7480 12784 7616
tri 12784 7480 12920 7616 nw
tri 10744 7344 10880 7480 sw
tri 10880 7344 11016 7480 se
rect 11016 7344 11424 7480
tri 11424 7344 11560 7480 sw
tri 11560 7344 11696 7480 se
rect 11696 7344 12104 7480
tri 12104 7344 12240 7480 sw
rect 10200 6936 12240 7344
tri 10200 6800 10336 6936 ne
rect 10336 6800 10744 6936
tri 10744 6800 10880 6936 nw
tri 10880 6800 11016 6936 ne
rect 11016 6800 11424 6936
tri 11424 6800 11560 6936 nw
tri 11560 6800 11696 6936 ne
rect 11696 6800 12104 6936
tri 12104 6800 12240 6936 nw
tri 13600 7344 13736 7480 se
rect 13736 7344 14144 7480
tri 14144 7344 14280 7480 sw
rect 13600 6936 14280 7344
tri 13600 6800 13736 6936 ne
rect 13736 6800 14144 6936
tri 14144 6800 14280 6936 nw
tri 9384 6664 9520 6800 sw
tri 9520 6664 9656 6800 se
rect 9656 6664 10064 6800
tri 10064 6664 10200 6800 sw
rect 7480 6256 10200 6664
tri 7480 6120 7616 6256 ne
tri 7480 5984 7616 6120 se
rect 7616 5984 8024 6256
tri 8024 6120 8160 6256 nw
tri 8160 6120 8296 6256 ne
tri 8024 5984 8160 6120 sw
tri 8160 5984 8296 6120 se
rect 8296 5984 8704 6256
tri 8704 6120 8840 6256 nw
tri 8840 6120 8976 6256 ne
rect 8976 6120 9384 6256
tri 9384 6120 9520 6256 nw
tri 9520 6120 9656 6256 ne
rect 9656 6120 10064 6256
tri 10064 6120 10200 6256 nw
tri 12920 6664 13056 6800 se
rect 13056 6664 13464 6800
tri 13464 6664 13600 6800 sw
rect 12920 6256 13600 6664
tri 12920 6120 13056 6256 ne
rect 13056 6120 13464 6256
tri 13464 6120 13600 6256 nw
tri 8704 5984 8840 6120 sw
rect 7480 5576 8840 5984
tri 7480 5440 7616 5576 ne
tri 5984 5304 6120 5440 sw
rect 5440 4896 6120 5304
tri 5440 4760 5576 4896 ne
tri 0 4624 136 4760 se
rect 136 4624 544 4760
tri 544 4624 680 4760 sw
tri 680 4624 816 4760 se
rect 816 4624 1224 4760
tri 1224 4624 1360 4760 sw
tri 1360 4624 1496 4760 se
rect 1496 4624 1904 4760
tri 1904 4624 2040 4760 sw
tri 2040 4624 2176 4760 se
rect 2176 4624 2584 4760
tri 2584 4624 2720 4760 sw
tri 2720 4624 2856 4760 se
rect 2856 4624 3264 4760
tri 3264 4624 3400 4760 sw
tri 3400 4624 3536 4760 se
rect 3536 4624 3944 4760
tri 3944 4624 4080 4760 sw
tri 4080 4624 4216 4760 se
rect 4216 4624 4624 4760
tri 4624 4624 4760 4760 sw
rect 0 4216 4760 4624
tri 0 4080 136 4216 ne
tri 0 3944 136 4080 se
rect 136 3944 544 4216
tri 544 4080 680 4216 nw
tri 680 4080 816 4216 ne
rect 816 4080 1224 4216
tri 1224 4080 1360 4216 nw
tri 1360 4080 1496 4216 ne
rect 1496 4080 1904 4216
tri 1904 4080 2040 4216 nw
tri 2040 4080 2176 4216 ne
rect 2176 4080 2584 4216
tri 2584 4080 2720 4216 nw
tri 2720 4080 2856 4216 ne
rect 2856 4080 3264 4216
tri 3264 4080 3400 4216 nw
tri 3400 4080 3536 4216 ne
rect 3536 4080 3944 4216
tri 3944 4080 4080 4216 nw
tri 4080 4080 4216 4216 ne
tri 544 3944 680 4080 sw
rect 0 3536 680 3944
tri 0 3400 136 3536 ne
tri 0 3264 136 3400 se
rect 136 3264 544 3536
tri 544 3400 680 3536 nw
tri 4080 3944 4216 4080 se
rect 4216 3944 4624 4216
tri 4624 4080 4760 4216 nw
tri 5440 4624 5576 4760 se
rect 5576 4624 5984 4896
tri 5984 4760 6120 4896 nw
tri 6800 5304 6936 5440 se
rect 6936 5304 7344 5440
tri 7344 5304 7480 5440 sw
tri 7480 5304 7616 5440 se
rect 7616 5304 8024 5576
tri 8024 5440 8160 5576 nw
tri 8160 5440 8296 5576 ne
tri 8024 5304 8160 5440 sw
tri 8160 5304 8296 5440 se
rect 8296 5304 8704 5576
tri 8704 5440 8840 5576 nw
tri 10880 5984 11016 6120 se
rect 11016 5984 11424 6120
tri 11424 5984 11560 6120 sw
rect 10880 5576 11560 5984
tri 10880 5440 11016 5576 ne
rect 11016 5440 11424 5576
tri 11424 5440 11560 5576 nw
tri 12240 5984 12376 6120 se
rect 12376 5984 12784 6120
tri 12784 5984 12920 6120 sw
rect 12240 5576 12920 5984
tri 12240 5440 12376 5576 ne
rect 12376 5440 12784 5576
tri 12784 5440 12920 5576 nw
tri 8704 5304 8840 5440 sw
tri 8840 5304 8976 5440 se
rect 8976 5304 9384 5440
tri 9384 5304 9520 5440 sw
rect 6800 4896 9520 5304
tri 6800 4760 6936 4896 ne
tri 5984 4624 6120 4760 sw
tri 6120 4624 6256 4760 se
rect 6256 4624 6664 4760
tri 6664 4624 6800 4760 sw
tri 6800 4624 6936 4760 se
rect 6936 4624 7344 4896
tri 7344 4760 7480 4896 nw
tri 7480 4760 7616 4896 ne
tri 7344 4624 7480 4760 sw
tri 7480 4624 7616 4760 se
rect 7616 4624 8024 4896
tri 8024 4760 8160 4896 nw
tri 8160 4760 8296 4896 ne
tri 8024 4624 8160 4760 sw
tri 8160 4624 8296 4760 se
rect 8296 4624 8704 4896
tri 8704 4760 8840 4896 nw
tri 8840 4760 8976 4896 ne
rect 8976 4760 9384 4896
tri 9384 4760 9520 4896 nw
tri 10200 5304 10336 5440 se
rect 10336 5304 10744 5440
tri 10744 5304 10880 5440 sw
rect 10200 4896 10880 5304
tri 10200 4760 10336 4896 ne
rect 10336 4760 10744 4896
tri 10744 4760 10880 4896 nw
tri 11560 5304 11696 5440 se
rect 11696 5304 12104 5440
tri 12104 5304 12240 5440 sw
rect 11560 4896 12240 5304
tri 11560 4760 11696 4896 ne
rect 11696 4760 12104 4896
tri 12104 4760 12240 4896 nw
tri 13600 5304 13736 5440 se
rect 13736 5304 14144 5440
tri 14144 5304 14280 5440 sw
rect 13600 4896 14280 5304
tri 13600 4760 13736 4896 ne
rect 13736 4760 14144 4896
tri 14144 4760 14280 4896 nw
tri 8704 4624 8840 4760 sw
rect 5440 4216 8840 4624
tri 5440 4080 5576 4216 ne
rect 5576 4080 5984 4216
tri 5984 4080 6120 4216 nw
tri 6120 4080 6256 4216 ne
rect 6256 4080 6664 4216
tri 6664 4080 6800 4216 nw
tri 6800 4080 6936 4216 ne
rect 6936 4080 7344 4216
tri 7344 4080 7480 4216 nw
tri 7480 4080 7616 4216 ne
rect 7616 4080 8024 4216
tri 8024 4080 8160 4216 nw
tri 8160 4080 8296 4216 ne
rect 8296 4080 8704 4216
tri 8704 4080 8840 4216 nw
tri 10880 4624 11016 4760 se
rect 11016 4624 11424 4760
tri 11424 4624 11560 4760 sw
rect 10880 4216 11560 4624
tri 10880 4080 11016 4216 ne
rect 11016 4080 11424 4216
tri 11424 4080 11560 4216 nw
tri 12920 4624 13056 4760 se
rect 13056 4624 13464 4760
tri 13464 4624 13600 4760 sw
rect 12920 4216 13600 4624
tri 12920 4080 13056 4216 ne
rect 13056 4080 13464 4216
tri 13464 4080 13600 4216 nw
tri 4624 3944 4760 4080 sw
rect 4080 3536 4760 3944
tri 4080 3400 4216 3536 ne
tri 544 3264 680 3400 sw
rect 0 2856 680 3264
tri 0 2720 136 2856 ne
tri 0 2584 136 2720 se
rect 136 2584 544 2856
tri 544 2720 680 2856 nw
tri 544 2584 680 2720 sw
rect 0 2176 680 2584
tri 0 2040 136 2176 ne
tri 0 1904 136 2040 se
rect 136 1904 544 2176
tri 544 2040 680 2176 nw
tri 544 1904 680 2040 sw
rect 0 1496 680 1904
tri 0 1360 136 1496 ne
tri 0 1224 136 1360 se
rect 136 1224 544 1496
tri 544 1360 680 1496 nw
tri 1360 3264 1496 3400 se
rect 1496 3264 1904 3400
tri 1904 3264 2040 3400 sw
tri 2040 3264 2176 3400 se
rect 2176 3264 2584 3400
tri 2584 3264 2720 3400 sw
tri 2720 3264 2856 3400 se
rect 2856 3264 3264 3400
tri 3264 3264 3400 3400 sw
rect 1360 2856 3400 3264
tri 1360 2720 1496 2856 ne
tri 1360 2584 1496 2720 se
rect 1496 2584 1904 2856
tri 1904 2720 2040 2856 nw
tri 2040 2720 2176 2856 ne
tri 1904 2584 2040 2720 sw
tri 2040 2584 2176 2720 se
rect 2176 2584 2584 2856
tri 2584 2720 2720 2856 nw
tri 2720 2720 2856 2856 ne
tri 2584 2584 2720 2720 sw
tri 2720 2584 2856 2720 se
rect 2856 2584 3264 2856
tri 3264 2720 3400 2856 nw
tri 3264 2584 3400 2720 sw
rect 1360 2176 3400 2584
tri 1360 2040 1496 2176 ne
tri 1360 1904 1496 2040 se
rect 1496 1904 1904 2176
tri 1904 2040 2040 2176 nw
tri 2040 2040 2176 2176 ne
tri 1904 1904 2040 2040 sw
tri 2040 1904 2176 2040 se
rect 2176 1904 2584 2176
tri 2584 2040 2720 2176 nw
tri 2720 2040 2856 2176 ne
tri 2584 1904 2720 2040 sw
tri 2720 1904 2856 2040 se
rect 2856 1904 3264 2176
tri 3264 2040 3400 2176 nw
tri 3264 1904 3400 2040 sw
rect 1360 1496 3400 1904
tri 1360 1360 1496 1496 ne
rect 1496 1360 1904 1496
tri 1904 1360 2040 1496 nw
tri 2040 1360 2176 1496 ne
rect 2176 1360 2584 1496
tri 2584 1360 2720 1496 nw
tri 2720 1360 2856 1496 ne
rect 2856 1360 3264 1496
tri 3264 1360 3400 1496 nw
tri 4080 3264 4216 3400 se
rect 4216 3264 4624 3536
tri 4624 3400 4760 3536 nw
tri 9520 3944 9656 4080 se
rect 9656 3944 10064 4080
tri 10064 3944 10200 4080 sw
rect 9520 3536 10200 3944
tri 9520 3400 9656 3536 ne
tri 4624 3264 4760 3400 sw
rect 4080 2856 4760 3264
tri 4080 2720 4216 2856 ne
tri 4080 2584 4216 2720 se
rect 4216 2584 4624 2856
tri 4624 2720 4760 2856 nw
tri 6120 3264 6256 3400 se
rect 6256 3264 6664 3400
tri 6664 3264 6800 3400 sw
tri 6800 3264 6936 3400 se
rect 6936 3264 7344 3400
tri 7344 3264 7480 3400 sw
tri 7480 3264 7616 3400 se
rect 7616 3264 8024 3400
tri 8024 3264 8160 3400 sw
rect 6120 2856 8160 3264
tri 6120 2720 6256 2856 ne
rect 6256 2720 6664 2856
tri 6664 2720 6800 2856 nw
tri 6800 2720 6936 2856 ne
tri 4624 2584 4760 2720 sw
rect 4080 2176 4760 2584
tri 4080 2040 4216 2176 ne
tri 4080 1904 4216 2040 se
rect 4216 1904 4624 2176
tri 4624 2040 4760 2176 nw
tri 4624 1904 4760 2040 sw
rect 4080 1496 4760 1904
tri 4080 1360 4216 1496 ne
tri 544 1224 680 1360 sw
rect 0 816 680 1224
tri 0 680 136 816 ne
tri 0 544 136 680 se
rect 136 544 544 816
tri 544 680 680 816 nw
tri 4080 1224 4216 1360 se
rect 4216 1224 4624 1496
tri 4624 1360 4760 1496 nw
tri 5440 2584 5576 2720 se
rect 5576 2584 5984 2720
tri 5984 2584 6120 2720 sw
rect 5440 2176 6120 2584
tri 5440 2040 5576 2176 ne
tri 5440 1904 5576 2040 se
rect 5576 1904 5984 2176
tri 5984 2040 6120 2176 nw
tri 6800 2584 6936 2720 se
rect 6936 2584 7344 2856
tri 7344 2720 7480 2856 nw
tri 7480 2720 7616 2856 ne
rect 7616 2720 8024 2856
tri 8024 2720 8160 2856 nw
tri 9520 3264 9656 3400 se
rect 9656 3264 10064 3536
tri 10064 3400 10200 3536 nw
tri 12240 3944 12376 4080 se
rect 12376 3944 12784 4080
tri 12784 3944 12920 4080 sw
rect 12240 3536 12920 3944
tri 12240 3400 12376 3536 ne
rect 12376 3400 12784 3536
tri 12784 3400 12920 3536 nw
tri 13600 3944 13736 4080 se
rect 13736 3944 14144 4080
tri 14144 3944 14280 4080 sw
rect 13600 3536 14280 3944
tri 13600 3400 13736 3536 ne
tri 10064 3264 10200 3400 sw
rect 9520 2856 10200 3264
tri 9520 2720 9656 2856 ne
tri 7344 2584 7480 2720 sw
rect 6800 2176 7480 2584
tri 6800 2040 6936 2176 ne
rect 6936 2040 7344 2176
tri 7344 2040 7480 2176 nw
tri 8160 2584 8296 2720 se
rect 8296 2584 8704 2720
tri 8704 2584 8840 2720 sw
rect 8160 2176 8840 2584
tri 8160 2040 8296 2176 ne
rect 8296 2040 8704 2176
tri 8704 2040 8840 2176 nw
tri 9520 2584 9656 2720 se
rect 9656 2584 10064 2856
tri 10064 2720 10200 2856 nw
tri 11560 3264 11696 3400 se
rect 11696 3264 12104 3400
tri 12104 3264 12240 3400 sw
rect 11560 2856 12240 3264
tri 11560 2720 11696 2856 ne
rect 11696 2720 12104 2856
tri 12104 2720 12240 2856 nw
tri 13600 3264 13736 3400 se
rect 13736 3264 14144 3536
tri 14144 3400 14280 3536 nw
tri 14144 3264 14280 3400 sw
rect 13600 2856 14280 3264
tri 13600 2720 13736 2856 ne
rect 13736 2720 14144 2856
tri 14144 2720 14280 2856 nw
tri 10064 2584 10200 2720 sw
rect 9520 2176 10200 2584
tri 9520 2040 9656 2176 ne
rect 9656 2040 10064 2176
tri 10064 2040 10200 2176 nw
tri 10880 2584 11016 2720 se
rect 11016 2584 11424 2720
tri 11424 2584 11560 2720 sw
rect 10880 2176 11560 2584
tri 10880 2040 11016 2176 ne
tri 5984 1904 6120 2040 sw
rect 5440 1496 6120 1904
tri 5440 1360 5576 1496 ne
rect 5576 1360 5984 1496
tri 5984 1360 6120 1496 nw
tri 7480 1904 7616 2040 se
rect 7616 1904 8024 2040
tri 8024 1904 8160 2040 sw
rect 7480 1496 8160 1904
tri 7480 1360 7616 1496 ne
tri 4624 1224 4760 1360 sw
rect 4080 816 4760 1224
tri 4080 680 4216 816 ne
tri 544 544 680 680 sw
tri 680 544 816 680 se
rect 816 544 1224 680
tri 1224 544 1360 680 sw
tri 1360 544 1496 680 se
rect 1496 544 1904 680
tri 1904 544 2040 680 sw
tri 2040 544 2176 680 se
rect 2176 544 2584 680
tri 2584 544 2720 680 sw
tri 2720 544 2856 680 se
rect 2856 544 3264 680
tri 3264 544 3400 680 sw
tri 3400 544 3536 680 se
rect 3536 544 3944 680
tri 3944 544 4080 680 sw
tri 4080 544 4216 680 se
rect 4216 544 4624 816
tri 4624 680 4760 816 nw
tri 6120 1224 6256 1360 se
rect 6256 1224 6664 1360
tri 6664 1224 6800 1360 sw
tri 6800 1224 6936 1360 se
rect 6936 1224 7344 1360
tri 7344 1224 7480 1360 sw
tri 7480 1224 7616 1360 se
rect 7616 1224 8024 1496
tri 8024 1360 8160 1496 nw
tri 10880 1904 11016 2040 se
rect 11016 1904 11424 2176
tri 11424 2040 11560 2176 nw
tri 12920 2584 13056 2720 se
rect 13056 2584 13464 2720
tri 13464 2584 13600 2720 sw
rect 12920 2176 13600 2584
tri 12920 2040 13056 2176 ne
rect 13056 2040 13464 2176
tri 13464 2040 13600 2176 nw
tri 11424 1904 11560 2040 sw
rect 10880 1496 11560 1904
tri 10880 1360 11016 1496 ne
tri 8024 1224 8160 1360 sw
rect 6120 816 8160 1224
tri 6120 680 6256 816 ne
rect 6256 680 6664 816
tri 6664 680 6800 816 nw
tri 6800 680 6936 816 ne
rect 6936 680 7344 816
tri 7344 680 7480 816 nw
tri 7480 680 7616 816 ne
rect 7616 680 8024 816
tri 8024 680 8160 816 nw
tri 8840 1224 8976 1360 se
rect 8976 1224 9384 1360
tri 9384 1224 9520 1360 sw
rect 8840 816 9520 1224
tri 8840 680 8976 816 ne
rect 8976 680 9384 816
tri 9384 680 9520 816 nw
tri 10880 1224 11016 1360 se
rect 11016 1224 11424 1496
tri 11424 1360 11560 1496 nw
tri 12240 1904 12376 2040 se
rect 12376 1904 12784 2040
tri 12784 1904 12920 2040 sw
rect 12240 1496 12920 1904
tri 12240 1360 12376 1496 ne
rect 12376 1360 12784 1496
tri 12784 1360 12920 1496 nw
tri 11424 1224 11560 1360 sw
tri 11560 1224 11696 1360 se
rect 11696 1224 12104 1360
tri 12104 1224 12240 1360 sw
rect 10880 816 12240 1224
tri 10880 680 11016 816 ne
rect 11016 680 11424 816
tri 11424 680 11560 816 nw
tri 11560 680 11696 816 ne
rect 11696 680 12104 816
tri 12104 680 12240 816 nw
tri 12920 1224 13056 1360 se
rect 13056 1224 13464 1360
tri 13464 1224 13600 1360 sw
tri 13600 1224 13736 1360 se
rect 13736 1224 14144 1360
tri 14144 1224 14280 1360 sw
rect 12920 816 14280 1224
tri 12920 680 13056 816 ne
tri 4624 544 4760 680 sw
rect 0 136 4760 544
tri 0 0 136 136 ne
rect 136 0 544 136
tri 544 0 680 136 nw
tri 680 0 816 136 ne
rect 816 0 1224 136
tri 1224 0 1360 136 nw
tri 1360 0 1496 136 ne
rect 1496 0 1904 136
tri 1904 0 2040 136 nw
tri 2040 0 2176 136 ne
rect 2176 0 2584 136
tri 2584 0 2720 136 nw
tri 2720 0 2856 136 ne
rect 2856 0 3264 136
tri 3264 0 3400 136 nw
tri 3400 0 3536 136 ne
rect 3536 0 3944 136
tri 3944 0 4080 136 nw
tri 4080 0 4216 136 ne
rect 4216 0 4624 136
tri 4624 0 4760 136 nw
tri 8160 544 8296 680 se
rect 8296 544 8704 680
tri 8704 544 8840 680 sw
rect 8160 136 8840 544
tri 8160 0 8296 136 ne
rect 8296 0 8704 136
tri 8704 0 8840 136 nw
tri 10200 544 10336 680 se
rect 10336 544 10744 680
tri 10744 544 10880 680 sw
rect 10200 136 10880 544
tri 10200 0 10336 136 ne
rect 10336 0 10744 136
tri 10744 0 10880 136 nw
tri 12920 544 13056 680 se
rect 13056 544 13464 816
tri 13464 680 13600 816 nw
tri 13600 680 13736 816 ne
rect 13736 680 14144 816
tri 14144 680 14280 816 nw
tri 13464 544 13600 680 sw
rect 12920 136 13600 544
tri 12920 0 13056 136 ne
rect 13056 0 13464 136
tri 13464 0 13600 136 nw
<< metal5 >>
tri 0 14144 136 14280 se
rect 136 14144 544 14280
tri 544 14144 680 14280 sw
tri 680 14144 816 14280 se
rect 816 14144 1224 14280
tri 1224 14144 1360 14280 sw
tri 1360 14144 1496 14280 se
rect 1496 14144 1904 14280
tri 1904 14144 2040 14280 sw
tri 2040 14144 2176 14280 se
rect 2176 14144 2584 14280
tri 2584 14144 2720 14280 sw
tri 2720 14144 2856 14280 se
rect 2856 14144 3264 14280
tri 3264 14144 3400 14280 sw
tri 3400 14144 3536 14280 se
rect 3536 14144 3944 14280
tri 3944 14144 4080 14280 sw
tri 4080 14144 4216 14280 se
rect 4216 14144 4624 14280
tri 4624 14144 4760 14280 sw
rect 0 13736 4760 14144
tri 0 13600 136 13736 ne
tri 0 13464 136 13600 se
rect 136 13464 544 13736
tri 544 13600 680 13736 nw
tri 680 13600 816 13736 ne
rect 816 13600 1224 13736
tri 1224 13600 1360 13736 nw
tri 1360 13600 1496 13736 ne
rect 1496 13600 1904 13736
tri 1904 13600 2040 13736 nw
tri 2040 13600 2176 13736 ne
rect 2176 13600 2584 13736
tri 2584 13600 2720 13736 nw
tri 2720 13600 2856 13736 ne
rect 2856 13600 3264 13736
tri 3264 13600 3400 13736 nw
tri 3400 13600 3536 13736 ne
rect 3536 13600 3944 13736
tri 3944 13600 4080 13736 nw
tri 4080 13600 4216 13736 ne
tri 544 13464 680 13600 sw
rect 0 13056 680 13464
tri 0 12920 136 13056 ne
tri 0 12784 136 12920 se
rect 136 12784 544 13056
tri 544 12920 680 13056 nw
tri 4080 13464 4216 13600 se
rect 4216 13464 4624 13736
tri 4624 13600 4760 13736 nw
tri 6120 14144 6256 14280 se
rect 6256 14144 6664 14280
tri 6664 14144 6800 14280 sw
tri 6800 14144 6936 14280 se
rect 6936 14144 7344 14280
tri 7344 14144 7480 14280 sw
rect 6120 13736 7480 14144
tri 6120 13600 6256 13736 ne
rect 6256 13600 6664 13736
tri 6664 13600 6800 13736 nw
tri 6800 13600 6936 13736 ne
tri 4624 13464 4760 13600 sw
rect 4080 13056 4760 13464
tri 4080 12920 4216 13056 ne
tri 544 12784 680 12920 sw
rect 0 12376 680 12784
tri 0 12240 136 12376 ne
tri 0 12104 136 12240 se
rect 136 12104 544 12376
tri 544 12240 680 12376 nw
tri 544 12104 680 12240 sw
rect 0 11696 680 12104
tri 0 11560 136 11696 ne
tri 0 11424 136 11560 se
rect 136 11424 544 11696
tri 544 11560 680 11696 nw
tri 544 11424 680 11560 sw
rect 0 11016 680 11424
tri 0 10880 136 11016 ne
tri 0 10744 136 10880 se
rect 136 10744 544 11016
tri 544 10880 680 11016 nw
tri 1360 12784 1496 12920 se
rect 1496 12784 1904 12920
tri 1904 12784 2040 12920 sw
tri 2040 12784 2176 12920 se
rect 2176 12784 2584 12920
tri 2584 12784 2720 12920 sw
tri 2720 12784 2856 12920 se
rect 2856 12784 3264 12920
tri 3264 12784 3400 12920 sw
rect 1360 12376 3400 12784
tri 1360 12240 1496 12376 ne
tri 1360 12104 1496 12240 se
rect 1496 12104 1904 12376
tri 1904 12240 2040 12376 nw
tri 2040 12240 2176 12376 ne
tri 1904 12104 2040 12240 sw
tri 2040 12104 2176 12240 se
rect 2176 12104 2584 12376
tri 2584 12240 2720 12376 nw
tri 2720 12240 2856 12376 ne
tri 2584 12104 2720 12240 sw
tri 2720 12104 2856 12240 se
rect 2856 12104 3264 12376
tri 3264 12240 3400 12376 nw
tri 3264 12104 3400 12240 sw
rect 1360 11696 3400 12104
tri 1360 11560 1496 11696 ne
tri 1360 11424 1496 11560 se
rect 1496 11424 1904 11696
tri 1904 11560 2040 11696 nw
tri 2040 11560 2176 11696 ne
tri 1904 11424 2040 11560 sw
tri 2040 11424 2176 11560 se
rect 2176 11424 2584 11696
tri 2584 11560 2720 11696 nw
tri 2720 11560 2856 11696 ne
tri 2584 11424 2720 11560 sw
tri 2720 11424 2856 11560 se
rect 2856 11424 3264 11696
tri 3264 11560 3400 11696 nw
tri 3264 11424 3400 11560 sw
rect 1360 11016 3400 11424
tri 1360 10880 1496 11016 ne
rect 1496 10880 1904 11016
tri 1904 10880 2040 11016 nw
tri 2040 10880 2176 11016 ne
rect 2176 10880 2584 11016
tri 2584 10880 2720 11016 nw
tri 2720 10880 2856 11016 ne
rect 2856 10880 3264 11016
tri 3264 10880 3400 11016 nw
tri 4080 12784 4216 12920 se
rect 4216 12784 4624 13056
tri 4624 12920 4760 13056 nw
tri 6800 13464 6936 13600 se
rect 6936 13464 7344 13736
tri 7344 13600 7480 13736 nw
tri 8160 14144 8296 14280 se
rect 8296 14144 8704 14280
tri 8704 14144 8840 14280 sw
rect 8160 13736 8840 14144
tri 8160 13600 8296 13736 ne
rect 8296 13600 8704 13736
tri 8704 13600 8840 13736 nw
tri 9520 14144 9656 14280 se
rect 9656 14144 10064 14280
tri 10064 14144 10200 14280 sw
tri 10200 14144 10336 14280 se
rect 10336 14144 10744 14280
tri 10744 14144 10880 14280 sw
tri 10880 14144 11016 14280 se
rect 11016 14144 11424 14280
tri 11424 14144 11560 14280 sw
tri 11560 14144 11696 14280 se
rect 11696 14144 12104 14280
tri 12104 14144 12240 14280 sw
tri 12240 14144 12376 14280 se
rect 12376 14144 12784 14280
tri 12784 14144 12920 14280 sw
tri 12920 14144 13056 14280 se
rect 13056 14144 13464 14280
tri 13464 14144 13600 14280 sw
tri 13600 14144 13736 14280 se
rect 13736 14144 14144 14280
tri 14144 14144 14280 14280 sw
rect 9520 13736 14280 14144
tri 9520 13600 9656 13736 ne
tri 7344 13464 7480 13600 sw
tri 7480 13464 7616 13600 se
rect 7616 13464 8024 13600
tri 8024 13464 8160 13600 sw
rect 6800 13056 8160 13464
tri 6800 12920 6936 13056 ne
rect 6936 12920 7344 13056
tri 7344 12920 7480 13056 nw
tri 7480 12920 7616 13056 ne
tri 4624 12784 4760 12920 sw
rect 4080 12376 4760 12784
tri 4080 12240 4216 12376 ne
tri 4080 12104 4216 12240 se
rect 4216 12104 4624 12376
tri 4624 12240 4760 12376 nw
tri 7480 12784 7616 12920 se
rect 7616 12784 8024 13056
tri 8024 12920 8160 13056 nw
tri 9520 13464 9656 13600 se
rect 9656 13464 10064 13736
tri 10064 13600 10200 13736 nw
tri 10200 13600 10336 13736 ne
rect 10336 13600 10744 13736
tri 10744 13600 10880 13736 nw
tri 10880 13600 11016 13736 ne
rect 11016 13600 11424 13736
tri 11424 13600 11560 13736 nw
tri 11560 13600 11696 13736 ne
rect 11696 13600 12104 13736
tri 12104 13600 12240 13736 nw
tri 12240 13600 12376 13736 ne
rect 12376 13600 12784 13736
tri 12784 13600 12920 13736 nw
tri 12920 13600 13056 13736 ne
rect 13056 13600 13464 13736
tri 13464 13600 13600 13736 nw
tri 13600 13600 13736 13736 ne
tri 10064 13464 10200 13600 sw
rect 9520 13056 10200 13464
tri 9520 12920 9656 13056 ne
tri 8024 12784 8160 12920 sw
tri 8160 12784 8296 12920 se
rect 8296 12784 8704 12920
tri 8704 12784 8840 12920 sw
rect 7480 12376 8840 12784
tri 7480 12240 7616 12376 ne
tri 4624 12104 4760 12240 sw
rect 4080 11696 4760 12104
tri 4080 11560 4216 11696 ne
tri 4080 11424 4216 11560 se
rect 4216 11424 4624 11696
tri 4624 11560 4760 11696 nw
tri 6120 12104 6256 12240 se
rect 6256 12104 6664 12240
tri 6664 12104 6800 12240 sw
rect 6120 11696 6800 12104
tri 6120 11560 6256 11696 ne
tri 4624 11424 4760 11560 sw
rect 4080 11016 4760 11424
tri 4080 10880 4216 11016 ne
tri 544 10744 680 10880 sw
rect 0 10336 680 10744
tri 0 10200 136 10336 ne
tri 0 10064 136 10200 se
rect 136 10064 544 10336
tri 544 10200 680 10336 nw
tri 4080 10744 4216 10880 se
rect 4216 10744 4624 11016
tri 4624 10880 4760 11016 nw
tri 5440 11424 5576 11560 se
rect 5576 11424 5984 11560
tri 5984 11424 6120 11560 sw
tri 6120 11424 6256 11560 se
rect 6256 11424 6664 11696
tri 6664 11560 6800 11696 nw
tri 7480 12104 7616 12240 se
rect 7616 12104 8024 12376
tri 8024 12240 8160 12376 nw
tri 8160 12240 8296 12376 ne
tri 8024 12104 8160 12240 sw
tri 8160 12104 8296 12240 se
rect 8296 12104 8704 12376
tri 8704 12240 8840 12376 nw
tri 8704 12104 8840 12240 sw
rect 7480 11696 8840 12104
tri 7480 11560 7616 11696 ne
rect 7616 11560 8024 11696
tri 8024 11560 8160 11696 nw
tri 8160 11560 8296 11696 ne
rect 8296 11560 8704 11696
tri 8704 11560 8840 11696 nw
tri 9520 12784 9656 12920 se
rect 9656 12784 10064 13056
tri 10064 12920 10200 13056 nw
tri 13600 13464 13736 13600 se
rect 13736 13464 14144 13736
tri 14144 13600 14280 13736 nw
tri 14144 13464 14280 13600 sw
rect 13600 13056 14280 13464
tri 13600 12920 13736 13056 ne
tri 10064 12784 10200 12920 sw
rect 9520 12376 10200 12784
tri 9520 12240 9656 12376 ne
tri 9520 12104 9656 12240 se
rect 9656 12104 10064 12376
tri 10064 12240 10200 12376 nw
tri 10064 12104 10200 12240 sw
rect 9520 11696 10200 12104
tri 9520 11560 9656 11696 ne
tri 6664 11424 6800 11560 sw
rect 5440 11016 6800 11424
tri 5440 10880 5576 11016 ne
rect 5576 10880 5984 11016
tri 5984 10880 6120 11016 nw
tri 6120 10880 6256 11016 ne
tri 4624 10744 4760 10880 sw
rect 4080 10336 4760 10744
tri 4080 10200 4216 10336 ne
tri 544 10064 680 10200 sw
tri 680 10064 816 10200 se
rect 816 10064 1224 10200
tri 1224 10064 1360 10200 sw
tri 1360 10064 1496 10200 se
rect 1496 10064 1904 10200
tri 1904 10064 2040 10200 sw
tri 2040 10064 2176 10200 se
rect 2176 10064 2584 10200
tri 2584 10064 2720 10200 sw
tri 2720 10064 2856 10200 se
rect 2856 10064 3264 10200
tri 3264 10064 3400 10200 sw
tri 3400 10064 3536 10200 se
rect 3536 10064 3944 10200
tri 3944 10064 4080 10200 sw
tri 4080 10064 4216 10200 se
rect 4216 10064 4624 10336
tri 4624 10200 4760 10336 nw
tri 6120 10744 6256 10880 se
rect 6256 10744 6664 11016
tri 6664 10880 6800 11016 nw
tri 9520 11424 9656 11560 se
rect 9656 11424 10064 11696
tri 10064 11560 10200 11696 nw
tri 10064 11424 10200 11560 sw
rect 9520 11016 10200 11424
tri 9520 10880 9656 11016 ne
tri 6664 10744 6800 10880 sw
tri 6800 10744 6936 10880 se
rect 6936 10744 7344 10880
tri 7344 10744 7480 10880 sw
rect 6120 10336 7480 10744
tri 6120 10200 6256 10336 ne
rect 6256 10200 6664 10336
tri 6664 10200 6800 10336 nw
tri 6800 10200 6936 10336 ne
tri 4624 10064 4760 10200 sw
rect 0 9656 4760 10064
tri 0 9520 136 9656 ne
rect 136 9520 544 9656
tri 544 9520 680 9656 nw
tri 680 9520 816 9656 ne
rect 816 9520 1224 9656
tri 1224 9520 1360 9656 nw
tri 1360 9520 1496 9656 ne
rect 1496 9520 1904 9656
tri 1904 9520 2040 9656 nw
tri 2040 9520 2176 9656 ne
rect 2176 9520 2584 9656
tri 2584 9520 2720 9656 nw
tri 2720 9520 2856 9656 ne
rect 2856 9520 3264 9656
tri 3264 9520 3400 9656 nw
tri 3400 9520 3536 9656 ne
rect 3536 9520 3944 9656
tri 3944 9520 4080 9656 nw
tri 4080 9520 4216 9656 ne
rect 4216 9520 4624 9656
tri 4624 9520 4760 9656 nw
tri 5440 10064 5576 10200 se
rect 5576 10064 5984 10200
tri 5984 10064 6120 10200 sw
rect 5440 9656 6120 10064
tri 5440 9520 5576 9656 ne
tri 5440 9384 5576 9520 se
rect 5576 9384 5984 9656
tri 5984 9520 6120 9656 nw
tri 6800 10064 6936 10200 se
rect 6936 10064 7344 10336
tri 7344 10200 7480 10336 nw
tri 7344 10064 7480 10200 sw
rect 6800 9656 7480 10064
tri 6800 9520 6936 9656 ne
tri 5984 9384 6120 9520 sw
tri 6120 9384 6256 9520 se
rect 6256 9384 6664 9520
tri 6664 9384 6800 9520 sw
tri 6800 9384 6936 9520 se
rect 6936 9384 7344 9656
tri 7344 9520 7480 9656 nw
tri 8160 10744 8296 10880 se
rect 8296 10744 8704 10880
tri 8704 10744 8840 10880 sw
rect 8160 10336 8840 10744
tri 8160 10200 8296 10336 ne
tri 8160 10064 8296 10200 se
rect 8296 10064 8704 10336
tri 8704 10200 8840 10336 nw
tri 8704 10064 8840 10200 sw
rect 8160 9656 8840 10064
tri 8160 9520 8296 9656 ne
rect 8296 9520 8704 9656
tri 8704 9520 8840 9656 nw
tri 9520 10744 9656 10880 se
rect 9656 10744 10064 11016
tri 10064 10880 10200 11016 nw
tri 10880 12784 11016 12920 se
rect 11016 12784 11424 12920
tri 11424 12784 11560 12920 sw
tri 11560 12784 11696 12920 se
rect 11696 12784 12104 12920
tri 12104 12784 12240 12920 sw
tri 12240 12784 12376 12920 se
rect 12376 12784 12784 12920
tri 12784 12784 12920 12920 sw
rect 10880 12376 12920 12784
tri 10880 12240 11016 12376 ne
tri 10880 12104 11016 12240 se
rect 11016 12104 11424 12376
tri 11424 12240 11560 12376 nw
tri 11560 12240 11696 12376 ne
tri 11424 12104 11560 12240 sw
tri 11560 12104 11696 12240 se
rect 11696 12104 12104 12376
tri 12104 12240 12240 12376 nw
tri 12240 12240 12376 12376 ne
tri 12104 12104 12240 12240 sw
tri 12240 12104 12376 12240 se
rect 12376 12104 12784 12376
tri 12784 12240 12920 12376 nw
tri 12784 12104 12920 12240 sw
rect 10880 11696 12920 12104
tri 10880 11560 11016 11696 ne
tri 10880 11424 11016 11560 se
rect 11016 11424 11424 11696
tri 11424 11560 11560 11696 nw
tri 11560 11560 11696 11696 ne
tri 11424 11424 11560 11560 sw
tri 11560 11424 11696 11560 se
rect 11696 11424 12104 11696
tri 12104 11560 12240 11696 nw
tri 12240 11560 12376 11696 ne
tri 12104 11424 12240 11560 sw
tri 12240 11424 12376 11560 se
rect 12376 11424 12784 11696
tri 12784 11560 12920 11696 nw
tri 12784 11424 12920 11560 sw
rect 10880 11016 12920 11424
tri 10880 10880 11016 11016 ne
rect 11016 10880 11424 11016
tri 11424 10880 11560 11016 nw
tri 11560 10880 11696 11016 ne
rect 11696 10880 12104 11016
tri 12104 10880 12240 11016 nw
tri 12240 10880 12376 11016 ne
rect 12376 10880 12784 11016
tri 12784 10880 12920 11016 nw
tri 13600 12784 13736 12920 se
rect 13736 12784 14144 13056
tri 14144 12920 14280 13056 nw
tri 14144 12784 14280 12920 sw
rect 13600 12376 14280 12784
tri 13600 12240 13736 12376 ne
tri 13600 12104 13736 12240 se
rect 13736 12104 14144 12376
tri 14144 12240 14280 12376 nw
tri 14144 12104 14280 12240 sw
rect 13600 11696 14280 12104
tri 13600 11560 13736 11696 ne
tri 13600 11424 13736 11560 se
rect 13736 11424 14144 11696
tri 14144 11560 14280 11696 nw
tri 14144 11424 14280 11560 sw
rect 13600 11016 14280 11424
tri 13600 10880 13736 11016 ne
tri 10064 10744 10200 10880 sw
rect 9520 10336 10200 10744
tri 9520 10200 9656 10336 ne
tri 9520 10064 9656 10200 se
rect 9656 10064 10064 10336
tri 10064 10200 10200 10336 nw
tri 13600 10744 13736 10880 se
rect 13736 10744 14144 11016
tri 14144 10880 14280 11016 nw
tri 14144 10744 14280 10880 sw
rect 13600 10336 14280 10744
tri 13600 10200 13736 10336 ne
tri 10064 10064 10200 10200 sw
tri 10200 10064 10336 10200 se
rect 10336 10064 10744 10200
tri 10744 10064 10880 10200 sw
tri 10880 10064 11016 10200 se
rect 11016 10064 11424 10200
tri 11424 10064 11560 10200 sw
tri 11560 10064 11696 10200 se
rect 11696 10064 12104 10200
tri 12104 10064 12240 10200 sw
tri 12240 10064 12376 10200 se
rect 12376 10064 12784 10200
tri 12784 10064 12920 10200 sw
tri 12920 10064 13056 10200 se
rect 13056 10064 13464 10200
tri 13464 10064 13600 10200 sw
tri 13600 10064 13736 10200 se
rect 13736 10064 14144 10336
tri 14144 10200 14280 10336 nw
tri 14144 10064 14280 10200 sw
rect 9520 9656 14280 10064
tri 9520 9520 9656 9656 ne
rect 9656 9520 10064 9656
tri 10064 9520 10200 9656 nw
tri 10200 9520 10336 9656 ne
rect 10336 9520 10744 9656
tri 10744 9520 10880 9656 nw
tri 10880 9520 11016 9656 ne
rect 11016 9520 11424 9656
tri 11424 9520 11560 9656 nw
tri 11560 9520 11696 9656 ne
rect 11696 9520 12104 9656
tri 12104 9520 12240 9656 nw
tri 12240 9520 12376 9656 ne
rect 12376 9520 12784 9656
tri 12784 9520 12920 9656 nw
tri 12920 9520 13056 9656 ne
rect 13056 9520 13464 9656
tri 13464 9520 13600 9656 nw
tri 13600 9520 13736 9656 ne
rect 13736 9520 14144 9656
tri 14144 9520 14280 9656 nw
tri 7344 9384 7480 9520 sw
rect 5440 8976 7480 9384
tri 5440 8840 5576 8976 ne
tri 1360 8704 1496 8840 se
rect 1496 8704 1904 8840
tri 1904 8704 2040 8840 sw
tri 2040 8704 2176 8840 se
rect 2176 8704 2584 8840
tri 2584 8704 2720 8840 sw
rect 1360 8296 2720 8704
tri 1360 8160 1496 8296 ne
tri 1360 8024 1496 8160 se
rect 1496 8024 1904 8296
tri 1904 8160 2040 8296 nw
tri 2040 8160 2176 8296 ne
tri 1904 8024 2040 8160 sw
tri 2040 8024 2176 8160 se
rect 2176 8024 2584 8296
tri 2584 8160 2720 8296 nw
tri 4080 8704 4216 8840 se
rect 4216 8704 4624 8840
tri 4624 8704 4760 8840 sw
tri 4760 8704 4896 8840 se
rect 4896 8704 5304 8840
tri 5304 8704 5440 8840 sw
tri 5440 8704 5576 8840 se
rect 5576 8704 5984 8976
tri 5984 8840 6120 8976 nw
tri 6120 8840 6256 8976 ne
tri 5984 8704 6120 8840 sw
tri 6120 8704 6256 8840 se
rect 6256 8704 6664 8976
tri 6664 8840 6800 8976 nw
tri 6800 8840 6936 8976 ne
rect 6936 8840 7344 8976
tri 7344 8840 7480 8976 nw
tri 6664 8704 6800 8840 sw
rect 4080 8296 6800 8704
tri 4080 8160 4216 8296 ne
rect 4216 8160 4624 8296
tri 4624 8160 4760 8296 nw
tri 4760 8160 4896 8296 ne
tri 2584 8024 2720 8160 sw
rect 1360 7616 2720 8024
tri 1360 7480 1496 7616 ne
tri 0 7344 136 7480 se
rect 136 7344 544 7480
tri 544 7344 680 7480 sw
tri 680 7344 816 7480 se
rect 816 7344 1224 7480
tri 1224 7344 1360 7480 sw
tri 1360 7344 1496 7480 se
rect 1496 7344 1904 7616
tri 1904 7480 2040 7616 nw
tri 2040 7480 2176 7616 ne
tri 1904 7344 2040 7480 sw
tri 2040 7344 2176 7480 se
rect 2176 7344 2584 7616
tri 2584 7480 2720 7616 nw
tri 4760 8024 4896 8160 se
rect 4896 8024 5304 8296
tri 5304 8160 5440 8296 nw
tri 5440 8160 5576 8296 ne
tri 5304 8024 5440 8160 sw
tri 5440 8024 5576 8160 se
rect 5576 8024 5984 8296
tri 5984 8160 6120 8296 nw
tri 6120 8160 6256 8296 ne
tri 5984 8024 6120 8160 sw
tri 6120 8024 6256 8160 se
rect 6256 8024 6664 8296
tri 6664 8160 6800 8296 nw
tri 7480 8704 7616 8840 se
rect 7616 8704 8024 8840
tri 8024 8704 8160 8840 sw
rect 7480 8296 8160 8704
tri 7480 8160 7616 8296 ne
rect 7616 8160 8024 8296
tri 8024 8160 8160 8296 nw
tri 8840 8704 8976 8840 se
rect 8976 8704 9384 8840
tri 9384 8704 9520 8840 sw
tri 9520 8704 9656 8840 se
rect 9656 8704 10064 8840
tri 10064 8704 10200 8840 sw
rect 8840 8296 10200 8704
tri 8840 8160 8976 8296 ne
tri 6664 8024 6800 8160 sw
tri 6800 8024 6936 8160 se
rect 6936 8024 7344 8160
tri 7344 8024 7480 8160 sw
rect 4760 7616 7480 8024
tri 4760 7480 4896 7616 ne
tri 2584 7344 2720 7480 sw
tri 2720 7344 2856 7480 se
rect 2856 7344 3264 7480
tri 3264 7344 3400 7480 sw
tri 3400 7344 3536 7480 se
rect 3536 7344 3944 7480
tri 3944 7344 4080 7480 sw
tri 4080 7344 4216 7480 se
rect 4216 7344 4624 7480
tri 4624 7344 4760 7480 sw
tri 4760 7344 4896 7480 se
rect 4896 7344 5304 7616
tri 5304 7480 5440 7616 nw
tri 5440 7480 5576 7616 ne
rect 5576 7480 5984 7616
tri 5984 7480 6120 7616 nw
tri 6120 7480 6256 7616 ne
tri 5304 7344 5440 7480 sw
rect 0 6936 5440 7344
tri 0 6800 136 6936 ne
rect 136 6800 544 6936
tri 544 6800 680 6936 nw
tri 680 6800 816 6936 ne
tri 680 6664 816 6800 se
rect 816 6664 1224 6936
tri 1224 6800 1360 6936 nw
tri 1360 6800 1496 6936 ne
tri 1224 6664 1360 6800 sw
tri 1360 6664 1496 6800 se
rect 1496 6664 1904 6936
tri 1904 6800 2040 6936 nw
tri 2040 6800 2176 6936 ne
rect 2176 6800 2584 6936
tri 2584 6800 2720 6936 nw
tri 2720 6800 2856 6936 ne
tri 1904 6664 2040 6800 sw
rect 680 6256 2040 6664
tri 680 6120 816 6256 ne
rect 816 6120 1224 6256
tri 1224 6120 1360 6256 nw
tri 1360 6120 1496 6256 ne
rect 1496 6120 1904 6256
tri 1904 6120 2040 6256 nw
tri 2720 6664 2856 6800 se
rect 2856 6664 3264 6936
tri 3264 6800 3400 6936 nw
tri 3400 6800 3536 6936 ne
rect 3536 6800 3944 6936
tri 3944 6800 4080 6936 nw
tri 4080 6800 4216 6936 ne
rect 4216 6800 4624 6936
tri 4624 6800 4760 6936 nw
tri 4760 6800 4896 6936 ne
tri 3264 6664 3400 6800 sw
rect 2720 6256 3400 6664
tri 2720 6120 2856 6256 ne
tri 0 5984 136 6120 se
rect 136 5984 544 6120
tri 544 5984 680 6120 sw
rect 0 5576 680 5984
tri 0 5440 136 5576 ne
rect 136 5440 544 5576
tri 544 5440 680 5576 nw
tri 2720 5984 2856 6120 se
rect 2856 5984 3264 6256
tri 3264 6120 3400 6256 nw
tri 4760 6664 4896 6800 se
rect 4896 6664 5304 6936
tri 5304 6800 5440 6936 nw
tri 6120 7344 6256 7480 se
rect 6256 7344 6664 7616
tri 6664 7480 6800 7616 nw
tri 6800 7480 6936 7616 ne
rect 6936 7480 7344 7616
tri 7344 7480 7480 7616 nw
tri 8840 8024 8976 8160 se
rect 8976 8024 9384 8296
tri 9384 8160 9520 8296 nw
tri 9520 8160 9656 8296 ne
rect 9656 8160 10064 8296
tri 10064 8160 10200 8296 nw
tri 10880 8704 11016 8840 se
rect 11016 8704 11424 8840
tri 11424 8704 11560 8840 sw
rect 10880 8296 11560 8704
tri 10880 8160 11016 8296 ne
rect 11016 8160 11424 8296
tri 11424 8160 11560 8296 nw
tri 9384 8024 9520 8160 sw
rect 8840 7616 9520 8024
tri 8840 7480 8976 7616 ne
tri 6664 7344 6800 7480 sw
rect 6120 6936 6800 7344
tri 6120 6800 6256 6936 ne
tri 5304 6664 5440 6800 sw
tri 5440 6664 5576 6800 se
rect 5576 6664 5984 6800
tri 5984 6664 6120 6800 sw
tri 6120 6664 6256 6800 se
rect 6256 6664 6664 6936
tri 6664 6800 6800 6936 nw
tri 6664 6664 6800 6800 sw
rect 4760 6256 6800 6664
tri 4760 6120 4896 6256 ne
rect 4896 6120 5304 6256
tri 5304 6120 5440 6256 nw
tri 5440 6120 5576 6256 ne
tri 3264 5984 3400 6120 sw
tri 3400 5984 3536 6120 se
rect 3536 5984 3944 6120
tri 3944 5984 4080 6120 sw
tri 4080 5984 4216 6120 se
rect 4216 5984 4624 6120
tri 4624 5984 4760 6120 sw
rect 2720 5576 4760 5984
tri 2720 5440 2856 5576 ne
rect 2856 5440 3264 5576
tri 3264 5440 3400 5576 nw
tri 3400 5440 3536 5576 ne
rect 3536 5440 3944 5576
tri 3944 5440 4080 5576 nw
tri 4080 5440 4216 5576 ne
rect 4216 5440 4624 5576
tri 4624 5440 4760 5576 nw
tri 5440 5984 5576 6120 se
rect 5576 5984 5984 6256
tri 5984 6120 6120 6256 nw
tri 6120 6120 6256 6256 ne
tri 5984 5984 6120 6120 sw
tri 6120 5984 6256 6120 se
rect 6256 5984 6664 6256
tri 6664 6120 6800 6256 nw
tri 6664 5984 6800 6120 sw
rect 5440 5576 6800 5984
tri 5440 5440 5576 5576 ne
tri 5440 5304 5576 5440 se
rect 5576 5304 5984 5576
tri 5984 5440 6120 5576 nw
tri 6120 5440 6256 5576 ne
rect 6256 5440 6664 5576
tri 6664 5440 6800 5576 nw
tri 7480 7344 7616 7480 se
rect 7616 7344 8024 7480
tri 8024 7344 8160 7480 sw
rect 7480 6936 8160 7344
tri 7480 6800 7616 6936 ne
tri 7480 6664 7616 6800 se
rect 7616 6664 8024 6936
tri 8024 6800 8160 6936 nw
tri 8840 7344 8976 7480 se
rect 8976 7344 9384 7616
tri 9384 7480 9520 7616 nw
tri 9384 7344 9520 7480 sw
rect 8840 6936 9520 7344
tri 8840 6800 8976 6936 ne
tri 8024 6664 8160 6800 sw
tri 8160 6664 8296 6800 se
rect 8296 6664 8704 6800
tri 8704 6664 8840 6800 sw
tri 8840 6664 8976 6800 se
rect 8976 6664 9384 6936
tri 9384 6800 9520 6936 nw
tri 10200 8024 10336 8160 se
rect 10336 8024 10744 8160
tri 10744 8024 10880 8160 sw
rect 10200 7616 10880 8024
tri 10200 7480 10336 7616 ne
tri 10200 7344 10336 7480 se
rect 10336 7344 10744 7616
tri 10744 7480 10880 7616 nw
tri 12240 8024 12376 8160 se
rect 12376 8024 12784 8160
tri 12784 8024 12920 8160 sw
rect 12240 7616 12920 8024
tri 12240 7480 12376 7616 ne
rect 12376 7480 12784 7616
tri 12784 7480 12920 7616 nw
tri 10744 7344 10880 7480 sw
tri 10880 7344 11016 7480 se
rect 11016 7344 11424 7480
tri 11424 7344 11560 7480 sw
tri 11560 7344 11696 7480 se
rect 11696 7344 12104 7480
tri 12104 7344 12240 7480 sw
rect 10200 6936 12240 7344
tri 10200 6800 10336 6936 ne
rect 10336 6800 10744 6936
tri 10744 6800 10880 6936 nw
tri 10880 6800 11016 6936 ne
rect 11016 6800 11424 6936
tri 11424 6800 11560 6936 nw
tri 11560 6800 11696 6936 ne
rect 11696 6800 12104 6936
tri 12104 6800 12240 6936 nw
tri 13600 7344 13736 7480 se
rect 13736 7344 14144 7480
tri 14144 7344 14280 7480 sw
rect 13600 6936 14280 7344
tri 13600 6800 13736 6936 ne
rect 13736 6800 14144 6936
tri 14144 6800 14280 6936 nw
tri 9384 6664 9520 6800 sw
tri 9520 6664 9656 6800 se
rect 9656 6664 10064 6800
tri 10064 6664 10200 6800 sw
rect 7480 6256 10200 6664
tri 7480 6120 7616 6256 ne
tri 7480 5984 7616 6120 se
rect 7616 5984 8024 6256
tri 8024 6120 8160 6256 nw
tri 8160 6120 8296 6256 ne
tri 8024 5984 8160 6120 sw
tri 8160 5984 8296 6120 se
rect 8296 5984 8704 6256
tri 8704 6120 8840 6256 nw
tri 8840 6120 8976 6256 ne
rect 8976 6120 9384 6256
tri 9384 6120 9520 6256 nw
tri 9520 6120 9656 6256 ne
rect 9656 6120 10064 6256
tri 10064 6120 10200 6256 nw
tri 12920 6664 13056 6800 se
rect 13056 6664 13464 6800
tri 13464 6664 13600 6800 sw
rect 12920 6256 13600 6664
tri 12920 6120 13056 6256 ne
rect 13056 6120 13464 6256
tri 13464 6120 13600 6256 nw
tri 8704 5984 8840 6120 sw
rect 7480 5576 8840 5984
tri 7480 5440 7616 5576 ne
tri 5984 5304 6120 5440 sw
rect 5440 4896 6120 5304
tri 5440 4760 5576 4896 ne
tri 0 4624 136 4760 se
rect 136 4624 544 4760
tri 544 4624 680 4760 sw
tri 680 4624 816 4760 se
rect 816 4624 1224 4760
tri 1224 4624 1360 4760 sw
tri 1360 4624 1496 4760 se
rect 1496 4624 1904 4760
tri 1904 4624 2040 4760 sw
tri 2040 4624 2176 4760 se
rect 2176 4624 2584 4760
tri 2584 4624 2720 4760 sw
tri 2720 4624 2856 4760 se
rect 2856 4624 3264 4760
tri 3264 4624 3400 4760 sw
tri 3400 4624 3536 4760 se
rect 3536 4624 3944 4760
tri 3944 4624 4080 4760 sw
tri 4080 4624 4216 4760 se
rect 4216 4624 4624 4760
tri 4624 4624 4760 4760 sw
rect 0 4216 4760 4624
tri 0 4080 136 4216 ne
tri 0 3944 136 4080 se
rect 136 3944 544 4216
tri 544 4080 680 4216 nw
tri 680 4080 816 4216 ne
rect 816 4080 1224 4216
tri 1224 4080 1360 4216 nw
tri 1360 4080 1496 4216 ne
rect 1496 4080 1904 4216
tri 1904 4080 2040 4216 nw
tri 2040 4080 2176 4216 ne
rect 2176 4080 2584 4216
tri 2584 4080 2720 4216 nw
tri 2720 4080 2856 4216 ne
rect 2856 4080 3264 4216
tri 3264 4080 3400 4216 nw
tri 3400 4080 3536 4216 ne
rect 3536 4080 3944 4216
tri 3944 4080 4080 4216 nw
tri 4080 4080 4216 4216 ne
tri 544 3944 680 4080 sw
rect 0 3536 680 3944
tri 0 3400 136 3536 ne
tri 0 3264 136 3400 se
rect 136 3264 544 3536
tri 544 3400 680 3536 nw
tri 4080 3944 4216 4080 se
rect 4216 3944 4624 4216
tri 4624 4080 4760 4216 nw
tri 5440 4624 5576 4760 se
rect 5576 4624 5984 4896
tri 5984 4760 6120 4896 nw
tri 6800 5304 6936 5440 se
rect 6936 5304 7344 5440
tri 7344 5304 7480 5440 sw
tri 7480 5304 7616 5440 se
rect 7616 5304 8024 5576
tri 8024 5440 8160 5576 nw
tri 8160 5440 8296 5576 ne
tri 8024 5304 8160 5440 sw
tri 8160 5304 8296 5440 se
rect 8296 5304 8704 5576
tri 8704 5440 8840 5576 nw
tri 10880 5984 11016 6120 se
rect 11016 5984 11424 6120
tri 11424 5984 11560 6120 sw
rect 10880 5576 11560 5984
tri 10880 5440 11016 5576 ne
rect 11016 5440 11424 5576
tri 11424 5440 11560 5576 nw
tri 12240 5984 12376 6120 se
rect 12376 5984 12784 6120
tri 12784 5984 12920 6120 sw
rect 12240 5576 12920 5984
tri 12240 5440 12376 5576 ne
rect 12376 5440 12784 5576
tri 12784 5440 12920 5576 nw
tri 8704 5304 8840 5440 sw
tri 8840 5304 8976 5440 se
rect 8976 5304 9384 5440
tri 9384 5304 9520 5440 sw
rect 6800 4896 9520 5304
tri 6800 4760 6936 4896 ne
tri 5984 4624 6120 4760 sw
tri 6120 4624 6256 4760 se
rect 6256 4624 6664 4760
tri 6664 4624 6800 4760 sw
tri 6800 4624 6936 4760 se
rect 6936 4624 7344 4896
tri 7344 4760 7480 4896 nw
tri 7480 4760 7616 4896 ne
tri 7344 4624 7480 4760 sw
tri 7480 4624 7616 4760 se
rect 7616 4624 8024 4896
tri 8024 4760 8160 4896 nw
tri 8160 4760 8296 4896 ne
tri 8024 4624 8160 4760 sw
tri 8160 4624 8296 4760 se
rect 8296 4624 8704 4896
tri 8704 4760 8840 4896 nw
tri 8840 4760 8976 4896 ne
rect 8976 4760 9384 4896
tri 9384 4760 9520 4896 nw
tri 10200 5304 10336 5440 se
rect 10336 5304 10744 5440
tri 10744 5304 10880 5440 sw
rect 10200 4896 10880 5304
tri 10200 4760 10336 4896 ne
rect 10336 4760 10744 4896
tri 10744 4760 10880 4896 nw
tri 11560 5304 11696 5440 se
rect 11696 5304 12104 5440
tri 12104 5304 12240 5440 sw
rect 11560 4896 12240 5304
tri 11560 4760 11696 4896 ne
rect 11696 4760 12104 4896
tri 12104 4760 12240 4896 nw
tri 13600 5304 13736 5440 se
rect 13736 5304 14144 5440
tri 14144 5304 14280 5440 sw
rect 13600 4896 14280 5304
tri 13600 4760 13736 4896 ne
rect 13736 4760 14144 4896
tri 14144 4760 14280 4896 nw
tri 8704 4624 8840 4760 sw
rect 5440 4216 8840 4624
tri 5440 4080 5576 4216 ne
rect 5576 4080 5984 4216
tri 5984 4080 6120 4216 nw
tri 6120 4080 6256 4216 ne
rect 6256 4080 6664 4216
tri 6664 4080 6800 4216 nw
tri 6800 4080 6936 4216 ne
rect 6936 4080 7344 4216
tri 7344 4080 7480 4216 nw
tri 7480 4080 7616 4216 ne
rect 7616 4080 8024 4216
tri 8024 4080 8160 4216 nw
tri 8160 4080 8296 4216 ne
rect 8296 4080 8704 4216
tri 8704 4080 8840 4216 nw
tri 10880 4624 11016 4760 se
rect 11016 4624 11424 4760
tri 11424 4624 11560 4760 sw
rect 10880 4216 11560 4624
tri 10880 4080 11016 4216 ne
rect 11016 4080 11424 4216
tri 11424 4080 11560 4216 nw
tri 12920 4624 13056 4760 se
rect 13056 4624 13464 4760
tri 13464 4624 13600 4760 sw
rect 12920 4216 13600 4624
tri 12920 4080 13056 4216 ne
rect 13056 4080 13464 4216
tri 13464 4080 13600 4216 nw
tri 4624 3944 4760 4080 sw
rect 4080 3536 4760 3944
tri 4080 3400 4216 3536 ne
tri 544 3264 680 3400 sw
rect 0 2856 680 3264
tri 0 2720 136 2856 ne
tri 0 2584 136 2720 se
rect 136 2584 544 2856
tri 544 2720 680 2856 nw
tri 544 2584 680 2720 sw
rect 0 2176 680 2584
tri 0 2040 136 2176 ne
tri 0 1904 136 2040 se
rect 136 1904 544 2176
tri 544 2040 680 2176 nw
tri 544 1904 680 2040 sw
rect 0 1496 680 1904
tri 0 1360 136 1496 ne
tri 0 1224 136 1360 se
rect 136 1224 544 1496
tri 544 1360 680 1496 nw
tri 1360 3264 1496 3400 se
rect 1496 3264 1904 3400
tri 1904 3264 2040 3400 sw
tri 2040 3264 2176 3400 se
rect 2176 3264 2584 3400
tri 2584 3264 2720 3400 sw
tri 2720 3264 2856 3400 se
rect 2856 3264 3264 3400
tri 3264 3264 3400 3400 sw
rect 1360 2856 3400 3264
tri 1360 2720 1496 2856 ne
tri 1360 2584 1496 2720 se
rect 1496 2584 1904 2856
tri 1904 2720 2040 2856 nw
tri 2040 2720 2176 2856 ne
tri 1904 2584 2040 2720 sw
tri 2040 2584 2176 2720 se
rect 2176 2584 2584 2856
tri 2584 2720 2720 2856 nw
tri 2720 2720 2856 2856 ne
tri 2584 2584 2720 2720 sw
tri 2720 2584 2856 2720 se
rect 2856 2584 3264 2856
tri 3264 2720 3400 2856 nw
tri 3264 2584 3400 2720 sw
rect 1360 2176 3400 2584
tri 1360 2040 1496 2176 ne
tri 1360 1904 1496 2040 se
rect 1496 1904 1904 2176
tri 1904 2040 2040 2176 nw
tri 2040 2040 2176 2176 ne
tri 1904 1904 2040 2040 sw
tri 2040 1904 2176 2040 se
rect 2176 1904 2584 2176
tri 2584 2040 2720 2176 nw
tri 2720 2040 2856 2176 ne
tri 2584 1904 2720 2040 sw
tri 2720 1904 2856 2040 se
rect 2856 1904 3264 2176
tri 3264 2040 3400 2176 nw
tri 3264 1904 3400 2040 sw
rect 1360 1496 3400 1904
tri 1360 1360 1496 1496 ne
rect 1496 1360 1904 1496
tri 1904 1360 2040 1496 nw
tri 2040 1360 2176 1496 ne
rect 2176 1360 2584 1496
tri 2584 1360 2720 1496 nw
tri 2720 1360 2856 1496 ne
rect 2856 1360 3264 1496
tri 3264 1360 3400 1496 nw
tri 4080 3264 4216 3400 se
rect 4216 3264 4624 3536
tri 4624 3400 4760 3536 nw
tri 9520 3944 9656 4080 se
rect 9656 3944 10064 4080
tri 10064 3944 10200 4080 sw
rect 9520 3536 10200 3944
tri 9520 3400 9656 3536 ne
tri 4624 3264 4760 3400 sw
rect 4080 2856 4760 3264
tri 4080 2720 4216 2856 ne
tri 4080 2584 4216 2720 se
rect 4216 2584 4624 2856
tri 4624 2720 4760 2856 nw
tri 6120 3264 6256 3400 se
rect 6256 3264 6664 3400
tri 6664 3264 6800 3400 sw
tri 6800 3264 6936 3400 se
rect 6936 3264 7344 3400
tri 7344 3264 7480 3400 sw
tri 7480 3264 7616 3400 se
rect 7616 3264 8024 3400
tri 8024 3264 8160 3400 sw
rect 6120 2856 8160 3264
tri 6120 2720 6256 2856 ne
rect 6256 2720 6664 2856
tri 6664 2720 6800 2856 nw
tri 6800 2720 6936 2856 ne
tri 4624 2584 4760 2720 sw
rect 4080 2176 4760 2584
tri 4080 2040 4216 2176 ne
tri 4080 1904 4216 2040 se
rect 4216 1904 4624 2176
tri 4624 2040 4760 2176 nw
tri 4624 1904 4760 2040 sw
rect 4080 1496 4760 1904
tri 4080 1360 4216 1496 ne
tri 544 1224 680 1360 sw
rect 0 816 680 1224
tri 0 680 136 816 ne
tri 0 544 136 680 se
rect 136 544 544 816
tri 544 680 680 816 nw
tri 4080 1224 4216 1360 se
rect 4216 1224 4624 1496
tri 4624 1360 4760 1496 nw
tri 5440 2584 5576 2720 se
rect 5576 2584 5984 2720
tri 5984 2584 6120 2720 sw
rect 5440 2176 6120 2584
tri 5440 2040 5576 2176 ne
tri 5440 1904 5576 2040 se
rect 5576 1904 5984 2176
tri 5984 2040 6120 2176 nw
tri 6800 2584 6936 2720 se
rect 6936 2584 7344 2856
tri 7344 2720 7480 2856 nw
tri 7480 2720 7616 2856 ne
rect 7616 2720 8024 2856
tri 8024 2720 8160 2856 nw
tri 9520 3264 9656 3400 se
rect 9656 3264 10064 3536
tri 10064 3400 10200 3536 nw
tri 12240 3944 12376 4080 se
rect 12376 3944 12784 4080
tri 12784 3944 12920 4080 sw
rect 12240 3536 12920 3944
tri 12240 3400 12376 3536 ne
rect 12376 3400 12784 3536
tri 12784 3400 12920 3536 nw
tri 13600 3944 13736 4080 se
rect 13736 3944 14144 4080
tri 14144 3944 14280 4080 sw
rect 13600 3536 14280 3944
tri 13600 3400 13736 3536 ne
tri 10064 3264 10200 3400 sw
rect 9520 2856 10200 3264
tri 9520 2720 9656 2856 ne
tri 7344 2584 7480 2720 sw
rect 6800 2176 7480 2584
tri 6800 2040 6936 2176 ne
rect 6936 2040 7344 2176
tri 7344 2040 7480 2176 nw
tri 8160 2584 8296 2720 se
rect 8296 2584 8704 2720
tri 8704 2584 8840 2720 sw
rect 8160 2176 8840 2584
tri 8160 2040 8296 2176 ne
rect 8296 2040 8704 2176
tri 8704 2040 8840 2176 nw
tri 9520 2584 9656 2720 se
rect 9656 2584 10064 2856
tri 10064 2720 10200 2856 nw
tri 11560 3264 11696 3400 se
rect 11696 3264 12104 3400
tri 12104 3264 12240 3400 sw
rect 11560 2856 12240 3264
tri 11560 2720 11696 2856 ne
rect 11696 2720 12104 2856
tri 12104 2720 12240 2856 nw
tri 13600 3264 13736 3400 se
rect 13736 3264 14144 3536
tri 14144 3400 14280 3536 nw
tri 14144 3264 14280 3400 sw
rect 13600 2856 14280 3264
tri 13600 2720 13736 2856 ne
rect 13736 2720 14144 2856
tri 14144 2720 14280 2856 nw
tri 10064 2584 10200 2720 sw
rect 9520 2176 10200 2584
tri 9520 2040 9656 2176 ne
rect 9656 2040 10064 2176
tri 10064 2040 10200 2176 nw
tri 10880 2584 11016 2720 se
rect 11016 2584 11424 2720
tri 11424 2584 11560 2720 sw
rect 10880 2176 11560 2584
tri 10880 2040 11016 2176 ne
tri 5984 1904 6120 2040 sw
rect 5440 1496 6120 1904
tri 5440 1360 5576 1496 ne
rect 5576 1360 5984 1496
tri 5984 1360 6120 1496 nw
tri 7480 1904 7616 2040 se
rect 7616 1904 8024 2040
tri 8024 1904 8160 2040 sw
rect 7480 1496 8160 1904
tri 7480 1360 7616 1496 ne
tri 4624 1224 4760 1360 sw
rect 4080 816 4760 1224
tri 4080 680 4216 816 ne
tri 544 544 680 680 sw
tri 680 544 816 680 se
rect 816 544 1224 680
tri 1224 544 1360 680 sw
tri 1360 544 1496 680 se
rect 1496 544 1904 680
tri 1904 544 2040 680 sw
tri 2040 544 2176 680 se
rect 2176 544 2584 680
tri 2584 544 2720 680 sw
tri 2720 544 2856 680 se
rect 2856 544 3264 680
tri 3264 544 3400 680 sw
tri 3400 544 3536 680 se
rect 3536 544 3944 680
tri 3944 544 4080 680 sw
tri 4080 544 4216 680 se
rect 4216 544 4624 816
tri 4624 680 4760 816 nw
tri 6120 1224 6256 1360 se
rect 6256 1224 6664 1360
tri 6664 1224 6800 1360 sw
tri 6800 1224 6936 1360 se
rect 6936 1224 7344 1360
tri 7344 1224 7480 1360 sw
tri 7480 1224 7616 1360 se
rect 7616 1224 8024 1496
tri 8024 1360 8160 1496 nw
tri 10880 1904 11016 2040 se
rect 11016 1904 11424 2176
tri 11424 2040 11560 2176 nw
tri 12920 2584 13056 2720 se
rect 13056 2584 13464 2720
tri 13464 2584 13600 2720 sw
rect 12920 2176 13600 2584
tri 12920 2040 13056 2176 ne
rect 13056 2040 13464 2176
tri 13464 2040 13600 2176 nw
tri 11424 1904 11560 2040 sw
rect 10880 1496 11560 1904
tri 10880 1360 11016 1496 ne
tri 8024 1224 8160 1360 sw
rect 6120 816 8160 1224
tri 6120 680 6256 816 ne
rect 6256 680 6664 816
tri 6664 680 6800 816 nw
tri 6800 680 6936 816 ne
rect 6936 680 7344 816
tri 7344 680 7480 816 nw
tri 7480 680 7616 816 ne
rect 7616 680 8024 816
tri 8024 680 8160 816 nw
tri 8840 1224 8976 1360 se
rect 8976 1224 9384 1360
tri 9384 1224 9520 1360 sw
rect 8840 816 9520 1224
tri 8840 680 8976 816 ne
rect 8976 680 9384 816
tri 9384 680 9520 816 nw
tri 10880 1224 11016 1360 se
rect 11016 1224 11424 1496
tri 11424 1360 11560 1496 nw
tri 12240 1904 12376 2040 se
rect 12376 1904 12784 2040
tri 12784 1904 12920 2040 sw
rect 12240 1496 12920 1904
tri 12240 1360 12376 1496 ne
rect 12376 1360 12784 1496
tri 12784 1360 12920 1496 nw
tri 11424 1224 11560 1360 sw
tri 11560 1224 11696 1360 se
rect 11696 1224 12104 1360
tri 12104 1224 12240 1360 sw
rect 10880 816 12240 1224
tri 10880 680 11016 816 ne
rect 11016 680 11424 816
tri 11424 680 11560 816 nw
tri 11560 680 11696 816 ne
rect 11696 680 12104 816
tri 12104 680 12240 816 nw
tri 12920 1224 13056 1360 se
rect 13056 1224 13464 1360
tri 13464 1224 13600 1360 sw
tri 13600 1224 13736 1360 se
rect 13736 1224 14144 1360
tri 14144 1224 14280 1360 sw
rect 12920 816 14280 1224
tri 12920 680 13056 816 ne
tri 4624 544 4760 680 sw
rect 0 136 4760 544
tri 0 0 136 136 ne
rect 136 0 544 136
tri 544 0 680 136 nw
tri 680 0 816 136 ne
rect 816 0 1224 136
tri 1224 0 1360 136 nw
tri 1360 0 1496 136 ne
rect 1496 0 1904 136
tri 1904 0 2040 136 nw
tri 2040 0 2176 136 ne
rect 2176 0 2584 136
tri 2584 0 2720 136 nw
tri 2720 0 2856 136 ne
rect 2856 0 3264 136
tri 3264 0 3400 136 nw
tri 3400 0 3536 136 ne
rect 3536 0 3944 136
tri 3944 0 4080 136 nw
tri 4080 0 4216 136 ne
rect 4216 0 4624 136
tri 4624 0 4760 136 nw
tri 8160 544 8296 680 se
rect 8296 544 8704 680
tri 8704 544 8840 680 sw
rect 8160 136 8840 544
tri 8160 0 8296 136 ne
rect 8296 0 8704 136
tri 8704 0 8840 136 nw
tri 10200 544 10336 680 se
rect 10336 544 10744 680
tri 10744 544 10880 680 sw
rect 10200 136 10880 544
tri 10200 0 10336 136 ne
rect 10336 0 10744 136
tri 10744 0 10880 136 nw
tri 12920 544 13056 680 se
rect 13056 544 13464 816
tri 13464 680 13600 816 nw
tri 13600 680 13736 816 ne
rect 13736 680 14144 816
tri 14144 680 14280 816 nw
tri 13464 544 13600 680 sw
rect 12920 136 13600 544
tri 12920 0 13056 136 ne
rect 13056 0 13464 136
tri 13464 0 13600 136 nw
<< fillblock >>
rect 0 0 14280 14280
<< properties >>
string FIXED_BBOX 0 0 14280 14280
string GDS_END 105844
string GDS_FILE ../../gds/gf180mcu_ws_ip__id.gds
string GDS_START 112
<< end >>
