magic
tech gf180mcuD
magscale 1 10
timestamp 1765934810
use gf180mcu_ocd_sram_test  gf180mcu_ocd_sram_test_0
timestamp 1765934810
transform 1 0 1 0 1 0
box 5200 5200 781200 501000
use gf180mcu_ws_ip__id  gf180mcu_ws_ip__id_0 wafer_space
timestamp 1765407047
transform 1 0 5201 0 1 5200
box 0 0 28560 28560
use gf180mcu_ws_ip__logo  gf180mcu_ws_ip__logo_0 wafer_space
timestamp 1765407047
transform 1 0 752551 0 1 472350
box 0 0 28650 28650
use sealring  sealring_0 wafer_space
timestamp 1765407464
transform 1 0 0 0 1 0
box 0 0 786400 506200
<< end >>
