magic
tech gf180mcuD
magscale 1 10
timestamp 1765059587
<< checkpaint >>
rect 89752 146428 90065 146528
<< metal2 >>
rect 89752 146522 90065 146528
rect 89752 146436 89764 146522
rect 90054 146436 90065 146522
rect 89752 146428 90065 146436
<< via2 >>
rect 89764 146436 90054 146522
<< metal3 >>
rect 89752 146522 90065 146528
rect 89752 146436 89764 146522
rect 90054 146436 90065 146522
rect 89752 146428 90065 146436
<< end >>
