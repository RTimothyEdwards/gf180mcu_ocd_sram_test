magic
tech gf180mcuD
magscale 1 10
timestamp 1765934810
<< metal3 >>
rect 104 69624 1916 69634
rect 104 69568 114 69624
rect 170 69568 238 69624
rect 294 69568 362 69624
rect 418 69568 486 69624
rect 542 69568 610 69624
rect 666 69568 734 69624
rect 790 69568 858 69624
rect 914 69568 982 69624
rect 1038 69568 1106 69624
rect 1162 69568 1230 69624
rect 1286 69568 1354 69624
rect 1410 69568 1478 69624
rect 1534 69568 1602 69624
rect 1658 69568 1726 69624
rect 1782 69568 1850 69624
rect 1906 69568 1916 69624
rect 104 69500 1916 69568
rect 104 69444 114 69500
rect 170 69444 238 69500
rect 294 69444 362 69500
rect 418 69444 486 69500
rect 542 69444 610 69500
rect 666 69444 734 69500
rect 790 69444 858 69500
rect 914 69444 982 69500
rect 1038 69444 1106 69500
rect 1162 69444 1230 69500
rect 1286 69444 1354 69500
rect 1410 69444 1478 69500
rect 1534 69444 1602 69500
rect 1658 69444 1726 69500
rect 1782 69444 1850 69500
rect 1906 69444 1916 69500
rect 104 69376 1916 69444
rect 104 69320 114 69376
rect 170 69320 238 69376
rect 294 69320 362 69376
rect 418 69320 486 69376
rect 542 69320 610 69376
rect 666 69320 734 69376
rect 790 69320 858 69376
rect 914 69320 982 69376
rect 1038 69320 1106 69376
rect 1162 69320 1230 69376
rect 1286 69320 1354 69376
rect 1410 69320 1478 69376
rect 1534 69320 1602 69376
rect 1658 69320 1726 69376
rect 1782 69320 1850 69376
rect 1906 69320 1916 69376
rect 104 69252 1916 69320
rect 104 69196 114 69252
rect 170 69196 238 69252
rect 294 69196 362 69252
rect 418 69196 486 69252
rect 542 69196 610 69252
rect 666 69196 734 69252
rect 790 69196 858 69252
rect 914 69196 982 69252
rect 1038 69196 1106 69252
rect 1162 69196 1230 69252
rect 1286 69196 1354 69252
rect 1410 69196 1478 69252
rect 1534 69196 1602 69252
rect 1658 69196 1726 69252
rect 1782 69196 1850 69252
rect 1906 69196 1916 69252
rect 104 69128 1916 69196
rect 104 69072 114 69128
rect 170 69072 238 69128
rect 294 69072 362 69128
rect 418 69072 486 69128
rect 542 69072 610 69128
rect 666 69072 734 69128
rect 790 69072 858 69128
rect 914 69072 982 69128
rect 1038 69072 1106 69128
rect 1162 69072 1230 69128
rect 1286 69072 1354 69128
rect 1410 69072 1478 69128
rect 1534 69072 1602 69128
rect 1658 69072 1726 69128
rect 1782 69072 1850 69128
rect 1906 69072 1916 69128
rect 104 69004 1916 69072
rect 104 68948 114 69004
rect 170 68948 238 69004
rect 294 68948 362 69004
rect 418 68948 486 69004
rect 542 68948 610 69004
rect 666 68948 734 69004
rect 790 68948 858 69004
rect 914 68948 982 69004
rect 1038 68948 1106 69004
rect 1162 68948 1230 69004
rect 1286 68948 1354 69004
rect 1410 68948 1478 69004
rect 1534 68948 1602 69004
rect 1658 68948 1726 69004
rect 1782 68948 1850 69004
rect 1906 68948 1916 69004
rect 104 68880 1916 68948
rect 104 68824 114 68880
rect 170 68824 238 68880
rect 294 68824 362 68880
rect 418 68824 486 68880
rect 542 68824 610 68880
rect 666 68824 734 68880
rect 790 68824 858 68880
rect 914 68824 982 68880
rect 1038 68824 1106 68880
rect 1162 68824 1230 68880
rect 1286 68824 1354 68880
rect 1410 68824 1478 68880
rect 1534 68824 1602 68880
rect 1658 68824 1726 68880
rect 1782 68824 1850 68880
rect 1906 68824 1916 68880
rect 104 68756 1916 68824
rect 104 68700 114 68756
rect 170 68700 238 68756
rect 294 68700 362 68756
rect 418 68700 486 68756
rect 542 68700 610 68756
rect 666 68700 734 68756
rect 790 68700 858 68756
rect 914 68700 982 68756
rect 1038 68700 1106 68756
rect 1162 68700 1230 68756
rect 1286 68700 1354 68756
rect 1410 68700 1478 68756
rect 1534 68700 1602 68756
rect 1658 68700 1726 68756
rect 1782 68700 1850 68756
rect 1906 68700 1916 68756
rect 104 68632 1916 68700
rect 104 68576 114 68632
rect 170 68576 238 68632
rect 294 68576 362 68632
rect 418 68576 486 68632
rect 542 68576 610 68632
rect 666 68576 734 68632
rect 790 68576 858 68632
rect 914 68576 982 68632
rect 1038 68576 1106 68632
rect 1162 68576 1230 68632
rect 1286 68576 1354 68632
rect 1410 68576 1478 68632
rect 1534 68576 1602 68632
rect 1658 68576 1726 68632
rect 1782 68576 1850 68632
rect 1906 68576 1916 68632
rect 104 68508 1916 68576
rect 104 68452 114 68508
rect 170 68452 238 68508
rect 294 68452 362 68508
rect 418 68452 486 68508
rect 542 68452 610 68508
rect 666 68452 734 68508
rect 790 68452 858 68508
rect 914 68452 982 68508
rect 1038 68452 1106 68508
rect 1162 68452 1230 68508
rect 1286 68452 1354 68508
rect 1410 68452 1478 68508
rect 1534 68452 1602 68508
rect 1658 68452 1726 68508
rect 1782 68452 1850 68508
rect 1906 68452 1916 68508
rect 104 68442 1916 68452
rect 104 68094 1916 68104
rect 104 68038 114 68094
rect 170 68038 238 68094
rect 294 68038 362 68094
rect 418 68038 486 68094
rect 542 68038 610 68094
rect 666 68038 734 68094
rect 790 68038 858 68094
rect 914 68038 982 68094
rect 1038 68038 1106 68094
rect 1162 68038 1230 68094
rect 1286 68038 1354 68094
rect 1410 68038 1478 68094
rect 1534 68038 1602 68094
rect 1658 68038 1726 68094
rect 1782 68038 1850 68094
rect 1906 68038 1916 68094
rect 104 67970 1916 68038
rect 104 67914 114 67970
rect 170 67914 238 67970
rect 294 67914 362 67970
rect 418 67914 486 67970
rect 542 67914 610 67970
rect 666 67914 734 67970
rect 790 67914 858 67970
rect 914 67914 982 67970
rect 1038 67914 1106 67970
rect 1162 67914 1230 67970
rect 1286 67914 1354 67970
rect 1410 67914 1478 67970
rect 1534 67914 1602 67970
rect 1658 67914 1726 67970
rect 1782 67914 1850 67970
rect 1906 67914 1916 67970
rect 104 67846 1916 67914
rect 104 67790 114 67846
rect 170 67790 238 67846
rect 294 67790 362 67846
rect 418 67790 486 67846
rect 542 67790 610 67846
rect 666 67790 734 67846
rect 790 67790 858 67846
rect 914 67790 982 67846
rect 1038 67790 1106 67846
rect 1162 67790 1230 67846
rect 1286 67790 1354 67846
rect 1410 67790 1478 67846
rect 1534 67790 1602 67846
rect 1658 67790 1726 67846
rect 1782 67790 1850 67846
rect 1906 67790 1916 67846
rect 104 67722 1916 67790
rect 104 67666 114 67722
rect 170 67666 238 67722
rect 294 67666 362 67722
rect 418 67666 486 67722
rect 542 67666 610 67722
rect 666 67666 734 67722
rect 790 67666 858 67722
rect 914 67666 982 67722
rect 1038 67666 1106 67722
rect 1162 67666 1230 67722
rect 1286 67666 1354 67722
rect 1410 67666 1478 67722
rect 1534 67666 1602 67722
rect 1658 67666 1726 67722
rect 1782 67666 1850 67722
rect 1906 67666 1916 67722
rect 104 67598 1916 67666
rect 104 67542 114 67598
rect 170 67542 238 67598
rect 294 67542 362 67598
rect 418 67542 486 67598
rect 542 67542 610 67598
rect 666 67542 734 67598
rect 790 67542 858 67598
rect 914 67542 982 67598
rect 1038 67542 1106 67598
rect 1162 67542 1230 67598
rect 1286 67542 1354 67598
rect 1410 67542 1478 67598
rect 1534 67542 1602 67598
rect 1658 67542 1726 67598
rect 1782 67542 1850 67598
rect 1906 67542 1916 67598
rect 104 67474 1916 67542
rect 104 67418 114 67474
rect 170 67418 238 67474
rect 294 67418 362 67474
rect 418 67418 486 67474
rect 542 67418 610 67474
rect 666 67418 734 67474
rect 790 67418 858 67474
rect 914 67418 982 67474
rect 1038 67418 1106 67474
rect 1162 67418 1230 67474
rect 1286 67418 1354 67474
rect 1410 67418 1478 67474
rect 1534 67418 1602 67474
rect 1658 67418 1726 67474
rect 1782 67418 1850 67474
rect 1906 67418 1916 67474
rect 104 67350 1916 67418
rect 104 67294 114 67350
rect 170 67294 238 67350
rect 294 67294 362 67350
rect 418 67294 486 67350
rect 542 67294 610 67350
rect 666 67294 734 67350
rect 790 67294 858 67350
rect 914 67294 982 67350
rect 1038 67294 1106 67350
rect 1162 67294 1230 67350
rect 1286 67294 1354 67350
rect 1410 67294 1478 67350
rect 1534 67294 1602 67350
rect 1658 67294 1726 67350
rect 1782 67294 1850 67350
rect 1906 67294 1916 67350
rect 104 67226 1916 67294
rect 104 67170 114 67226
rect 170 67170 238 67226
rect 294 67170 362 67226
rect 418 67170 486 67226
rect 542 67170 610 67226
rect 666 67170 734 67226
rect 790 67170 858 67226
rect 914 67170 982 67226
rect 1038 67170 1106 67226
rect 1162 67170 1230 67226
rect 1286 67170 1354 67226
rect 1410 67170 1478 67226
rect 1534 67170 1602 67226
rect 1658 67170 1726 67226
rect 1782 67170 1850 67226
rect 1906 67170 1916 67226
rect 104 67102 1916 67170
rect 104 67046 114 67102
rect 170 67046 238 67102
rect 294 67046 362 67102
rect 418 67046 486 67102
rect 542 67046 610 67102
rect 666 67046 734 67102
rect 790 67046 858 67102
rect 914 67046 982 67102
rect 1038 67046 1106 67102
rect 1162 67046 1230 67102
rect 1286 67046 1354 67102
rect 1410 67046 1478 67102
rect 1534 67046 1602 67102
rect 1658 67046 1726 67102
rect 1782 67046 1850 67102
rect 1906 67046 1916 67102
rect 104 66978 1916 67046
rect 104 66922 114 66978
rect 170 66922 238 66978
rect 294 66922 362 66978
rect 418 66922 486 66978
rect 542 66922 610 66978
rect 666 66922 734 66978
rect 790 66922 858 66978
rect 914 66922 982 66978
rect 1038 66922 1106 66978
rect 1162 66922 1230 66978
rect 1286 66922 1354 66978
rect 1410 66922 1478 66978
rect 1534 66922 1602 66978
rect 1658 66922 1726 66978
rect 1782 66922 1850 66978
rect 1906 66922 1916 66978
rect 104 66912 1916 66922
rect 104 66484 1916 66494
rect 104 66428 114 66484
rect 170 66428 238 66484
rect 294 66428 362 66484
rect 418 66428 486 66484
rect 542 66428 610 66484
rect 666 66428 734 66484
rect 790 66428 858 66484
rect 914 66428 982 66484
rect 1038 66428 1106 66484
rect 1162 66428 1230 66484
rect 1286 66428 1354 66484
rect 1410 66428 1478 66484
rect 1534 66428 1602 66484
rect 1658 66428 1726 66484
rect 1782 66428 1850 66484
rect 1906 66428 1916 66484
rect 104 66360 1916 66428
rect 104 66304 114 66360
rect 170 66304 238 66360
rect 294 66304 362 66360
rect 418 66304 486 66360
rect 542 66304 610 66360
rect 666 66304 734 66360
rect 790 66304 858 66360
rect 914 66304 982 66360
rect 1038 66304 1106 66360
rect 1162 66304 1230 66360
rect 1286 66304 1354 66360
rect 1410 66304 1478 66360
rect 1534 66304 1602 66360
rect 1658 66304 1726 66360
rect 1782 66304 1850 66360
rect 1906 66304 1916 66360
rect 104 66236 1916 66304
rect 104 66180 114 66236
rect 170 66180 238 66236
rect 294 66180 362 66236
rect 418 66180 486 66236
rect 542 66180 610 66236
rect 666 66180 734 66236
rect 790 66180 858 66236
rect 914 66180 982 66236
rect 1038 66180 1106 66236
rect 1162 66180 1230 66236
rect 1286 66180 1354 66236
rect 1410 66180 1478 66236
rect 1534 66180 1602 66236
rect 1658 66180 1726 66236
rect 1782 66180 1850 66236
rect 1906 66180 1916 66236
rect 104 66112 1916 66180
rect 104 66056 114 66112
rect 170 66056 238 66112
rect 294 66056 362 66112
rect 418 66056 486 66112
rect 542 66056 610 66112
rect 666 66056 734 66112
rect 790 66056 858 66112
rect 914 66056 982 66112
rect 1038 66056 1106 66112
rect 1162 66056 1230 66112
rect 1286 66056 1354 66112
rect 1410 66056 1478 66112
rect 1534 66056 1602 66112
rect 1658 66056 1726 66112
rect 1782 66056 1850 66112
rect 1906 66056 1916 66112
rect 104 65988 1916 66056
rect 104 65932 114 65988
rect 170 65932 238 65988
rect 294 65932 362 65988
rect 418 65932 486 65988
rect 542 65932 610 65988
rect 666 65932 734 65988
rect 790 65932 858 65988
rect 914 65932 982 65988
rect 1038 65932 1106 65988
rect 1162 65932 1230 65988
rect 1286 65932 1354 65988
rect 1410 65932 1478 65988
rect 1534 65932 1602 65988
rect 1658 65932 1726 65988
rect 1782 65932 1850 65988
rect 1906 65932 1916 65988
rect 104 65864 1916 65932
rect 104 65808 114 65864
rect 170 65808 238 65864
rect 294 65808 362 65864
rect 418 65808 486 65864
rect 542 65808 610 65864
rect 666 65808 734 65864
rect 790 65808 858 65864
rect 914 65808 982 65864
rect 1038 65808 1106 65864
rect 1162 65808 1230 65864
rect 1286 65808 1354 65864
rect 1410 65808 1478 65864
rect 1534 65808 1602 65864
rect 1658 65808 1726 65864
rect 1782 65808 1850 65864
rect 1906 65808 1916 65864
rect 104 65740 1916 65808
rect 104 65684 114 65740
rect 170 65684 238 65740
rect 294 65684 362 65740
rect 418 65684 486 65740
rect 542 65684 610 65740
rect 666 65684 734 65740
rect 790 65684 858 65740
rect 914 65684 982 65740
rect 1038 65684 1106 65740
rect 1162 65684 1230 65740
rect 1286 65684 1354 65740
rect 1410 65684 1478 65740
rect 1534 65684 1602 65740
rect 1658 65684 1726 65740
rect 1782 65684 1850 65740
rect 1906 65684 1916 65740
rect 104 65616 1916 65684
rect 104 65560 114 65616
rect 170 65560 238 65616
rect 294 65560 362 65616
rect 418 65560 486 65616
rect 542 65560 610 65616
rect 666 65560 734 65616
rect 790 65560 858 65616
rect 914 65560 982 65616
rect 1038 65560 1106 65616
rect 1162 65560 1230 65616
rect 1286 65560 1354 65616
rect 1410 65560 1478 65616
rect 1534 65560 1602 65616
rect 1658 65560 1726 65616
rect 1782 65560 1850 65616
rect 1906 65560 1916 65616
rect 104 65492 1916 65560
rect 104 65436 114 65492
rect 170 65436 238 65492
rect 294 65436 362 65492
rect 418 65436 486 65492
rect 542 65436 610 65492
rect 666 65436 734 65492
rect 790 65436 858 65492
rect 914 65436 982 65492
rect 1038 65436 1106 65492
rect 1162 65436 1230 65492
rect 1286 65436 1354 65492
rect 1410 65436 1478 65492
rect 1534 65436 1602 65492
rect 1658 65436 1726 65492
rect 1782 65436 1850 65492
rect 1906 65436 1916 65492
rect 104 65368 1916 65436
rect 104 65312 114 65368
rect 170 65312 238 65368
rect 294 65312 362 65368
rect 418 65312 486 65368
rect 542 65312 610 65368
rect 666 65312 734 65368
rect 790 65312 858 65368
rect 914 65312 982 65368
rect 1038 65312 1106 65368
rect 1162 65312 1230 65368
rect 1286 65312 1354 65368
rect 1410 65312 1478 65368
rect 1534 65312 1602 65368
rect 1658 65312 1726 65368
rect 1782 65312 1850 65368
rect 1906 65312 1916 65368
rect 104 65302 1916 65312
rect 104 64886 1916 64896
rect 104 64830 114 64886
rect 170 64830 238 64886
rect 294 64830 362 64886
rect 418 64830 486 64886
rect 542 64830 610 64886
rect 666 64830 734 64886
rect 790 64830 858 64886
rect 914 64830 982 64886
rect 1038 64830 1106 64886
rect 1162 64830 1230 64886
rect 1286 64830 1354 64886
rect 1410 64830 1478 64886
rect 1534 64830 1602 64886
rect 1658 64830 1726 64886
rect 1782 64830 1850 64886
rect 1906 64830 1916 64886
rect 104 64762 1916 64830
rect 104 64706 114 64762
rect 170 64706 238 64762
rect 294 64706 362 64762
rect 418 64706 486 64762
rect 542 64706 610 64762
rect 666 64706 734 64762
rect 790 64706 858 64762
rect 914 64706 982 64762
rect 1038 64706 1106 64762
rect 1162 64706 1230 64762
rect 1286 64706 1354 64762
rect 1410 64706 1478 64762
rect 1534 64706 1602 64762
rect 1658 64706 1726 64762
rect 1782 64706 1850 64762
rect 1906 64706 1916 64762
rect 104 64638 1916 64706
rect 104 64582 114 64638
rect 170 64582 238 64638
rect 294 64582 362 64638
rect 418 64582 486 64638
rect 542 64582 610 64638
rect 666 64582 734 64638
rect 790 64582 858 64638
rect 914 64582 982 64638
rect 1038 64582 1106 64638
rect 1162 64582 1230 64638
rect 1286 64582 1354 64638
rect 1410 64582 1478 64638
rect 1534 64582 1602 64638
rect 1658 64582 1726 64638
rect 1782 64582 1850 64638
rect 1906 64582 1916 64638
rect 104 64514 1916 64582
rect 104 64458 114 64514
rect 170 64458 238 64514
rect 294 64458 362 64514
rect 418 64458 486 64514
rect 542 64458 610 64514
rect 666 64458 734 64514
rect 790 64458 858 64514
rect 914 64458 982 64514
rect 1038 64458 1106 64514
rect 1162 64458 1230 64514
rect 1286 64458 1354 64514
rect 1410 64458 1478 64514
rect 1534 64458 1602 64514
rect 1658 64458 1726 64514
rect 1782 64458 1850 64514
rect 1906 64458 1916 64514
rect 104 64390 1916 64458
rect 104 64334 114 64390
rect 170 64334 238 64390
rect 294 64334 362 64390
rect 418 64334 486 64390
rect 542 64334 610 64390
rect 666 64334 734 64390
rect 790 64334 858 64390
rect 914 64334 982 64390
rect 1038 64334 1106 64390
rect 1162 64334 1230 64390
rect 1286 64334 1354 64390
rect 1410 64334 1478 64390
rect 1534 64334 1602 64390
rect 1658 64334 1726 64390
rect 1782 64334 1850 64390
rect 1906 64334 1916 64390
rect 104 64266 1916 64334
rect 104 64210 114 64266
rect 170 64210 238 64266
rect 294 64210 362 64266
rect 418 64210 486 64266
rect 542 64210 610 64266
rect 666 64210 734 64266
rect 790 64210 858 64266
rect 914 64210 982 64266
rect 1038 64210 1106 64266
rect 1162 64210 1230 64266
rect 1286 64210 1354 64266
rect 1410 64210 1478 64266
rect 1534 64210 1602 64266
rect 1658 64210 1726 64266
rect 1782 64210 1850 64266
rect 1906 64210 1916 64266
rect 104 64142 1916 64210
rect 104 64086 114 64142
rect 170 64086 238 64142
rect 294 64086 362 64142
rect 418 64086 486 64142
rect 542 64086 610 64142
rect 666 64086 734 64142
rect 790 64086 858 64142
rect 914 64086 982 64142
rect 1038 64086 1106 64142
rect 1162 64086 1230 64142
rect 1286 64086 1354 64142
rect 1410 64086 1478 64142
rect 1534 64086 1602 64142
rect 1658 64086 1726 64142
rect 1782 64086 1850 64142
rect 1906 64086 1916 64142
rect 104 64018 1916 64086
rect 104 63962 114 64018
rect 170 63962 238 64018
rect 294 63962 362 64018
rect 418 63962 486 64018
rect 542 63962 610 64018
rect 666 63962 734 64018
rect 790 63962 858 64018
rect 914 63962 982 64018
rect 1038 63962 1106 64018
rect 1162 63962 1230 64018
rect 1286 63962 1354 64018
rect 1410 63962 1478 64018
rect 1534 63962 1602 64018
rect 1658 63962 1726 64018
rect 1782 63962 1850 64018
rect 1906 63962 1916 64018
rect 104 63894 1916 63962
rect 104 63838 114 63894
rect 170 63838 238 63894
rect 294 63838 362 63894
rect 418 63838 486 63894
rect 542 63838 610 63894
rect 666 63838 734 63894
rect 790 63838 858 63894
rect 914 63838 982 63894
rect 1038 63838 1106 63894
rect 1162 63838 1230 63894
rect 1286 63838 1354 63894
rect 1410 63838 1478 63894
rect 1534 63838 1602 63894
rect 1658 63838 1726 63894
rect 1782 63838 1850 63894
rect 1906 63838 1916 63894
rect 104 63770 1916 63838
rect 104 63714 114 63770
rect 170 63714 238 63770
rect 294 63714 362 63770
rect 418 63714 486 63770
rect 542 63714 610 63770
rect 666 63714 734 63770
rect 790 63714 858 63770
rect 914 63714 982 63770
rect 1038 63714 1106 63770
rect 1162 63714 1230 63770
rect 1286 63714 1354 63770
rect 1410 63714 1478 63770
rect 1534 63714 1602 63770
rect 1658 63714 1726 63770
rect 1782 63714 1850 63770
rect 1906 63714 1916 63770
rect 104 63704 1916 63714
rect 104 63295 1916 63305
rect 104 63239 114 63295
rect 170 63239 238 63295
rect 294 63239 362 63295
rect 418 63239 486 63295
rect 542 63239 610 63295
rect 666 63239 734 63295
rect 790 63239 858 63295
rect 914 63239 982 63295
rect 1038 63239 1106 63295
rect 1162 63239 1230 63295
rect 1286 63239 1354 63295
rect 1410 63239 1478 63295
rect 1534 63239 1602 63295
rect 1658 63239 1726 63295
rect 1782 63239 1850 63295
rect 1906 63239 1916 63295
rect 104 63171 1916 63239
rect 104 63115 114 63171
rect 170 63115 238 63171
rect 294 63115 362 63171
rect 418 63115 486 63171
rect 542 63115 610 63171
rect 666 63115 734 63171
rect 790 63115 858 63171
rect 914 63115 982 63171
rect 1038 63115 1106 63171
rect 1162 63115 1230 63171
rect 1286 63115 1354 63171
rect 1410 63115 1478 63171
rect 1534 63115 1602 63171
rect 1658 63115 1726 63171
rect 1782 63115 1850 63171
rect 1906 63115 1916 63171
rect 104 63047 1916 63115
rect 104 62991 114 63047
rect 170 62991 238 63047
rect 294 62991 362 63047
rect 418 62991 486 63047
rect 542 62991 610 63047
rect 666 62991 734 63047
rect 790 62991 858 63047
rect 914 62991 982 63047
rect 1038 62991 1106 63047
rect 1162 62991 1230 63047
rect 1286 62991 1354 63047
rect 1410 62991 1478 63047
rect 1534 62991 1602 63047
rect 1658 62991 1726 63047
rect 1782 62991 1850 63047
rect 1906 62991 1916 63047
rect 104 62923 1916 62991
rect 104 62867 114 62923
rect 170 62867 238 62923
rect 294 62867 362 62923
rect 418 62867 486 62923
rect 542 62867 610 62923
rect 666 62867 734 62923
rect 790 62867 858 62923
rect 914 62867 982 62923
rect 1038 62867 1106 62923
rect 1162 62867 1230 62923
rect 1286 62867 1354 62923
rect 1410 62867 1478 62923
rect 1534 62867 1602 62923
rect 1658 62867 1726 62923
rect 1782 62867 1850 62923
rect 1906 62867 1916 62923
rect 104 62799 1916 62867
rect 104 62743 114 62799
rect 170 62743 238 62799
rect 294 62743 362 62799
rect 418 62743 486 62799
rect 542 62743 610 62799
rect 666 62743 734 62799
rect 790 62743 858 62799
rect 914 62743 982 62799
rect 1038 62743 1106 62799
rect 1162 62743 1230 62799
rect 1286 62743 1354 62799
rect 1410 62743 1478 62799
rect 1534 62743 1602 62799
rect 1658 62743 1726 62799
rect 1782 62743 1850 62799
rect 1906 62743 1916 62799
rect 104 62675 1916 62743
rect 104 62619 114 62675
rect 170 62619 238 62675
rect 294 62619 362 62675
rect 418 62619 486 62675
rect 542 62619 610 62675
rect 666 62619 734 62675
rect 790 62619 858 62675
rect 914 62619 982 62675
rect 1038 62619 1106 62675
rect 1162 62619 1230 62675
rect 1286 62619 1354 62675
rect 1410 62619 1478 62675
rect 1534 62619 1602 62675
rect 1658 62619 1726 62675
rect 1782 62619 1850 62675
rect 1906 62619 1916 62675
rect 104 62551 1916 62619
rect 104 62495 114 62551
rect 170 62495 238 62551
rect 294 62495 362 62551
rect 418 62495 486 62551
rect 542 62495 610 62551
rect 666 62495 734 62551
rect 790 62495 858 62551
rect 914 62495 982 62551
rect 1038 62495 1106 62551
rect 1162 62495 1230 62551
rect 1286 62495 1354 62551
rect 1410 62495 1478 62551
rect 1534 62495 1602 62551
rect 1658 62495 1726 62551
rect 1782 62495 1850 62551
rect 1906 62495 1916 62551
rect 104 62427 1916 62495
rect 104 62371 114 62427
rect 170 62371 238 62427
rect 294 62371 362 62427
rect 418 62371 486 62427
rect 542 62371 610 62427
rect 666 62371 734 62427
rect 790 62371 858 62427
rect 914 62371 982 62427
rect 1038 62371 1106 62427
rect 1162 62371 1230 62427
rect 1286 62371 1354 62427
rect 1410 62371 1478 62427
rect 1534 62371 1602 62427
rect 1658 62371 1726 62427
rect 1782 62371 1850 62427
rect 1906 62371 1916 62427
rect 104 62303 1916 62371
rect 104 62247 114 62303
rect 170 62247 238 62303
rect 294 62247 362 62303
rect 418 62247 486 62303
rect 542 62247 610 62303
rect 666 62247 734 62303
rect 790 62247 858 62303
rect 914 62247 982 62303
rect 1038 62247 1106 62303
rect 1162 62247 1230 62303
rect 1286 62247 1354 62303
rect 1410 62247 1478 62303
rect 1534 62247 1602 62303
rect 1658 62247 1726 62303
rect 1782 62247 1850 62303
rect 1906 62247 1916 62303
rect 104 62179 1916 62247
rect 104 62123 114 62179
rect 170 62123 238 62179
rect 294 62123 362 62179
rect 418 62123 486 62179
rect 542 62123 610 62179
rect 666 62123 734 62179
rect 790 62123 858 62179
rect 914 62123 982 62179
rect 1038 62123 1106 62179
rect 1162 62123 1230 62179
rect 1286 62123 1354 62179
rect 1410 62123 1478 62179
rect 1534 62123 1602 62179
rect 1658 62123 1726 62179
rect 1782 62123 1850 62179
rect 1906 62123 1916 62179
rect 104 62113 1916 62123
rect 104 61695 1916 61705
rect 104 61639 114 61695
rect 170 61639 238 61695
rect 294 61639 362 61695
rect 418 61639 486 61695
rect 542 61639 610 61695
rect 666 61639 734 61695
rect 790 61639 858 61695
rect 914 61639 982 61695
rect 1038 61639 1106 61695
rect 1162 61639 1230 61695
rect 1286 61639 1354 61695
rect 1410 61639 1478 61695
rect 1534 61639 1602 61695
rect 1658 61639 1726 61695
rect 1782 61639 1850 61695
rect 1906 61639 1916 61695
rect 104 61571 1916 61639
rect 104 61515 114 61571
rect 170 61515 238 61571
rect 294 61515 362 61571
rect 418 61515 486 61571
rect 542 61515 610 61571
rect 666 61515 734 61571
rect 790 61515 858 61571
rect 914 61515 982 61571
rect 1038 61515 1106 61571
rect 1162 61515 1230 61571
rect 1286 61515 1354 61571
rect 1410 61515 1478 61571
rect 1534 61515 1602 61571
rect 1658 61515 1726 61571
rect 1782 61515 1850 61571
rect 1906 61515 1916 61571
rect 104 61447 1916 61515
rect 104 61391 114 61447
rect 170 61391 238 61447
rect 294 61391 362 61447
rect 418 61391 486 61447
rect 542 61391 610 61447
rect 666 61391 734 61447
rect 790 61391 858 61447
rect 914 61391 982 61447
rect 1038 61391 1106 61447
rect 1162 61391 1230 61447
rect 1286 61391 1354 61447
rect 1410 61391 1478 61447
rect 1534 61391 1602 61447
rect 1658 61391 1726 61447
rect 1782 61391 1850 61447
rect 1906 61391 1916 61447
rect 104 61323 1916 61391
rect 104 61267 114 61323
rect 170 61267 238 61323
rect 294 61267 362 61323
rect 418 61267 486 61323
rect 542 61267 610 61323
rect 666 61267 734 61323
rect 790 61267 858 61323
rect 914 61267 982 61323
rect 1038 61267 1106 61323
rect 1162 61267 1230 61323
rect 1286 61267 1354 61323
rect 1410 61267 1478 61323
rect 1534 61267 1602 61323
rect 1658 61267 1726 61323
rect 1782 61267 1850 61323
rect 1906 61267 1916 61323
rect 104 61199 1916 61267
rect 104 61143 114 61199
rect 170 61143 238 61199
rect 294 61143 362 61199
rect 418 61143 486 61199
rect 542 61143 610 61199
rect 666 61143 734 61199
rect 790 61143 858 61199
rect 914 61143 982 61199
rect 1038 61143 1106 61199
rect 1162 61143 1230 61199
rect 1286 61143 1354 61199
rect 1410 61143 1478 61199
rect 1534 61143 1602 61199
rect 1658 61143 1726 61199
rect 1782 61143 1850 61199
rect 1906 61143 1916 61199
rect 104 61075 1916 61143
rect 104 61019 114 61075
rect 170 61019 238 61075
rect 294 61019 362 61075
rect 418 61019 486 61075
rect 542 61019 610 61075
rect 666 61019 734 61075
rect 790 61019 858 61075
rect 914 61019 982 61075
rect 1038 61019 1106 61075
rect 1162 61019 1230 61075
rect 1286 61019 1354 61075
rect 1410 61019 1478 61075
rect 1534 61019 1602 61075
rect 1658 61019 1726 61075
rect 1782 61019 1850 61075
rect 1906 61019 1916 61075
rect 104 60951 1916 61019
rect 104 60895 114 60951
rect 170 60895 238 60951
rect 294 60895 362 60951
rect 418 60895 486 60951
rect 542 60895 610 60951
rect 666 60895 734 60951
rect 790 60895 858 60951
rect 914 60895 982 60951
rect 1038 60895 1106 60951
rect 1162 60895 1230 60951
rect 1286 60895 1354 60951
rect 1410 60895 1478 60951
rect 1534 60895 1602 60951
rect 1658 60895 1726 60951
rect 1782 60895 1850 60951
rect 1906 60895 1916 60951
rect 104 60827 1916 60895
rect 104 60771 114 60827
rect 170 60771 238 60827
rect 294 60771 362 60827
rect 418 60771 486 60827
rect 542 60771 610 60827
rect 666 60771 734 60827
rect 790 60771 858 60827
rect 914 60771 982 60827
rect 1038 60771 1106 60827
rect 1162 60771 1230 60827
rect 1286 60771 1354 60827
rect 1410 60771 1478 60827
rect 1534 60771 1602 60827
rect 1658 60771 1726 60827
rect 1782 60771 1850 60827
rect 1906 60771 1916 60827
rect 104 60703 1916 60771
rect 104 60647 114 60703
rect 170 60647 238 60703
rect 294 60647 362 60703
rect 418 60647 486 60703
rect 542 60647 610 60703
rect 666 60647 734 60703
rect 790 60647 858 60703
rect 914 60647 982 60703
rect 1038 60647 1106 60703
rect 1162 60647 1230 60703
rect 1286 60647 1354 60703
rect 1410 60647 1478 60703
rect 1534 60647 1602 60703
rect 1658 60647 1726 60703
rect 1782 60647 1850 60703
rect 1906 60647 1916 60703
rect 104 60579 1916 60647
rect 104 60523 114 60579
rect 170 60523 238 60579
rect 294 60523 362 60579
rect 418 60523 486 60579
rect 542 60523 610 60579
rect 666 60523 734 60579
rect 790 60523 858 60579
rect 914 60523 982 60579
rect 1038 60523 1106 60579
rect 1162 60523 1230 60579
rect 1286 60523 1354 60579
rect 1410 60523 1478 60579
rect 1534 60523 1602 60579
rect 1658 60523 1726 60579
rect 1782 60523 1850 60579
rect 1906 60523 1916 60579
rect 104 60513 1916 60523
rect 104 60090 1916 60100
rect 104 60034 114 60090
rect 170 60034 238 60090
rect 294 60034 362 60090
rect 418 60034 486 60090
rect 542 60034 610 60090
rect 666 60034 734 60090
rect 790 60034 858 60090
rect 914 60034 982 60090
rect 1038 60034 1106 60090
rect 1162 60034 1230 60090
rect 1286 60034 1354 60090
rect 1410 60034 1478 60090
rect 1534 60034 1602 60090
rect 1658 60034 1726 60090
rect 1782 60034 1850 60090
rect 1906 60034 1916 60090
rect 104 59966 1916 60034
rect 104 59910 114 59966
rect 170 59910 238 59966
rect 294 59910 362 59966
rect 418 59910 486 59966
rect 542 59910 610 59966
rect 666 59910 734 59966
rect 790 59910 858 59966
rect 914 59910 982 59966
rect 1038 59910 1106 59966
rect 1162 59910 1230 59966
rect 1286 59910 1354 59966
rect 1410 59910 1478 59966
rect 1534 59910 1602 59966
rect 1658 59910 1726 59966
rect 1782 59910 1850 59966
rect 1906 59910 1916 59966
rect 104 59842 1916 59910
rect 104 59786 114 59842
rect 170 59786 238 59842
rect 294 59786 362 59842
rect 418 59786 486 59842
rect 542 59786 610 59842
rect 666 59786 734 59842
rect 790 59786 858 59842
rect 914 59786 982 59842
rect 1038 59786 1106 59842
rect 1162 59786 1230 59842
rect 1286 59786 1354 59842
rect 1410 59786 1478 59842
rect 1534 59786 1602 59842
rect 1658 59786 1726 59842
rect 1782 59786 1850 59842
rect 1906 59786 1916 59842
rect 104 59718 1916 59786
rect 104 59662 114 59718
rect 170 59662 238 59718
rect 294 59662 362 59718
rect 418 59662 486 59718
rect 542 59662 610 59718
rect 666 59662 734 59718
rect 790 59662 858 59718
rect 914 59662 982 59718
rect 1038 59662 1106 59718
rect 1162 59662 1230 59718
rect 1286 59662 1354 59718
rect 1410 59662 1478 59718
rect 1534 59662 1602 59718
rect 1658 59662 1726 59718
rect 1782 59662 1850 59718
rect 1906 59662 1916 59718
rect 104 59594 1916 59662
rect 104 59538 114 59594
rect 170 59538 238 59594
rect 294 59538 362 59594
rect 418 59538 486 59594
rect 542 59538 610 59594
rect 666 59538 734 59594
rect 790 59538 858 59594
rect 914 59538 982 59594
rect 1038 59538 1106 59594
rect 1162 59538 1230 59594
rect 1286 59538 1354 59594
rect 1410 59538 1478 59594
rect 1534 59538 1602 59594
rect 1658 59538 1726 59594
rect 1782 59538 1850 59594
rect 1906 59538 1916 59594
rect 104 59470 1916 59538
rect 104 59414 114 59470
rect 170 59414 238 59470
rect 294 59414 362 59470
rect 418 59414 486 59470
rect 542 59414 610 59470
rect 666 59414 734 59470
rect 790 59414 858 59470
rect 914 59414 982 59470
rect 1038 59414 1106 59470
rect 1162 59414 1230 59470
rect 1286 59414 1354 59470
rect 1410 59414 1478 59470
rect 1534 59414 1602 59470
rect 1658 59414 1726 59470
rect 1782 59414 1850 59470
rect 1906 59414 1916 59470
rect 104 59346 1916 59414
rect 104 59290 114 59346
rect 170 59290 238 59346
rect 294 59290 362 59346
rect 418 59290 486 59346
rect 542 59290 610 59346
rect 666 59290 734 59346
rect 790 59290 858 59346
rect 914 59290 982 59346
rect 1038 59290 1106 59346
rect 1162 59290 1230 59346
rect 1286 59290 1354 59346
rect 1410 59290 1478 59346
rect 1534 59290 1602 59346
rect 1658 59290 1726 59346
rect 1782 59290 1850 59346
rect 1906 59290 1916 59346
rect 104 59222 1916 59290
rect 104 59166 114 59222
rect 170 59166 238 59222
rect 294 59166 362 59222
rect 418 59166 486 59222
rect 542 59166 610 59222
rect 666 59166 734 59222
rect 790 59166 858 59222
rect 914 59166 982 59222
rect 1038 59166 1106 59222
rect 1162 59166 1230 59222
rect 1286 59166 1354 59222
rect 1410 59166 1478 59222
rect 1534 59166 1602 59222
rect 1658 59166 1726 59222
rect 1782 59166 1850 59222
rect 1906 59166 1916 59222
rect 104 59098 1916 59166
rect 104 59042 114 59098
rect 170 59042 238 59098
rect 294 59042 362 59098
rect 418 59042 486 59098
rect 542 59042 610 59098
rect 666 59042 734 59098
rect 790 59042 858 59098
rect 914 59042 982 59098
rect 1038 59042 1106 59098
rect 1162 59042 1230 59098
rect 1286 59042 1354 59098
rect 1410 59042 1478 59098
rect 1534 59042 1602 59098
rect 1658 59042 1726 59098
rect 1782 59042 1850 59098
rect 1906 59042 1916 59098
rect 104 58974 1916 59042
rect 104 58918 114 58974
rect 170 58918 238 58974
rect 294 58918 362 58974
rect 418 58918 486 58974
rect 542 58918 610 58974
rect 666 58918 734 58974
rect 790 58918 858 58974
rect 914 58918 982 58974
rect 1038 58918 1106 58974
rect 1162 58918 1230 58974
rect 1286 58918 1354 58974
rect 1410 58918 1478 58974
rect 1534 58918 1602 58974
rect 1658 58918 1726 58974
rect 1782 58918 1850 58974
rect 1906 58918 1916 58974
rect 104 58908 1916 58918
rect 104 58485 1916 58495
rect 104 58429 114 58485
rect 170 58429 238 58485
rect 294 58429 362 58485
rect 418 58429 486 58485
rect 542 58429 610 58485
rect 666 58429 734 58485
rect 790 58429 858 58485
rect 914 58429 982 58485
rect 1038 58429 1106 58485
rect 1162 58429 1230 58485
rect 1286 58429 1354 58485
rect 1410 58429 1478 58485
rect 1534 58429 1602 58485
rect 1658 58429 1726 58485
rect 1782 58429 1850 58485
rect 1906 58429 1916 58485
rect 104 58361 1916 58429
rect 104 58305 114 58361
rect 170 58305 238 58361
rect 294 58305 362 58361
rect 418 58305 486 58361
rect 542 58305 610 58361
rect 666 58305 734 58361
rect 790 58305 858 58361
rect 914 58305 982 58361
rect 1038 58305 1106 58361
rect 1162 58305 1230 58361
rect 1286 58305 1354 58361
rect 1410 58305 1478 58361
rect 1534 58305 1602 58361
rect 1658 58305 1726 58361
rect 1782 58305 1850 58361
rect 1906 58305 1916 58361
rect 104 58237 1916 58305
rect 104 58181 114 58237
rect 170 58181 238 58237
rect 294 58181 362 58237
rect 418 58181 486 58237
rect 542 58181 610 58237
rect 666 58181 734 58237
rect 790 58181 858 58237
rect 914 58181 982 58237
rect 1038 58181 1106 58237
rect 1162 58181 1230 58237
rect 1286 58181 1354 58237
rect 1410 58181 1478 58237
rect 1534 58181 1602 58237
rect 1658 58181 1726 58237
rect 1782 58181 1850 58237
rect 1906 58181 1916 58237
rect 104 58113 1916 58181
rect 104 58057 114 58113
rect 170 58057 238 58113
rect 294 58057 362 58113
rect 418 58057 486 58113
rect 542 58057 610 58113
rect 666 58057 734 58113
rect 790 58057 858 58113
rect 914 58057 982 58113
rect 1038 58057 1106 58113
rect 1162 58057 1230 58113
rect 1286 58057 1354 58113
rect 1410 58057 1478 58113
rect 1534 58057 1602 58113
rect 1658 58057 1726 58113
rect 1782 58057 1850 58113
rect 1906 58057 1916 58113
rect 104 57989 1916 58057
rect 104 57933 114 57989
rect 170 57933 238 57989
rect 294 57933 362 57989
rect 418 57933 486 57989
rect 542 57933 610 57989
rect 666 57933 734 57989
rect 790 57933 858 57989
rect 914 57933 982 57989
rect 1038 57933 1106 57989
rect 1162 57933 1230 57989
rect 1286 57933 1354 57989
rect 1410 57933 1478 57989
rect 1534 57933 1602 57989
rect 1658 57933 1726 57989
rect 1782 57933 1850 57989
rect 1906 57933 1916 57989
rect 104 57865 1916 57933
rect 104 57809 114 57865
rect 170 57809 238 57865
rect 294 57809 362 57865
rect 418 57809 486 57865
rect 542 57809 610 57865
rect 666 57809 734 57865
rect 790 57809 858 57865
rect 914 57809 982 57865
rect 1038 57809 1106 57865
rect 1162 57809 1230 57865
rect 1286 57809 1354 57865
rect 1410 57809 1478 57865
rect 1534 57809 1602 57865
rect 1658 57809 1726 57865
rect 1782 57809 1850 57865
rect 1906 57809 1916 57865
rect 104 57741 1916 57809
rect 104 57685 114 57741
rect 170 57685 238 57741
rect 294 57685 362 57741
rect 418 57685 486 57741
rect 542 57685 610 57741
rect 666 57685 734 57741
rect 790 57685 858 57741
rect 914 57685 982 57741
rect 1038 57685 1106 57741
rect 1162 57685 1230 57741
rect 1286 57685 1354 57741
rect 1410 57685 1478 57741
rect 1534 57685 1602 57741
rect 1658 57685 1726 57741
rect 1782 57685 1850 57741
rect 1906 57685 1916 57741
rect 104 57617 1916 57685
rect 104 57561 114 57617
rect 170 57561 238 57617
rect 294 57561 362 57617
rect 418 57561 486 57617
rect 542 57561 610 57617
rect 666 57561 734 57617
rect 790 57561 858 57617
rect 914 57561 982 57617
rect 1038 57561 1106 57617
rect 1162 57561 1230 57617
rect 1286 57561 1354 57617
rect 1410 57561 1478 57617
rect 1534 57561 1602 57617
rect 1658 57561 1726 57617
rect 1782 57561 1850 57617
rect 1906 57561 1916 57617
rect 104 57493 1916 57561
rect 104 57437 114 57493
rect 170 57437 238 57493
rect 294 57437 362 57493
rect 418 57437 486 57493
rect 542 57437 610 57493
rect 666 57437 734 57493
rect 790 57437 858 57493
rect 914 57437 982 57493
rect 1038 57437 1106 57493
rect 1162 57437 1230 57493
rect 1286 57437 1354 57493
rect 1410 57437 1478 57493
rect 1534 57437 1602 57493
rect 1658 57437 1726 57493
rect 1782 57437 1850 57493
rect 1906 57437 1916 57493
rect 104 57369 1916 57437
rect 104 57313 114 57369
rect 170 57313 238 57369
rect 294 57313 362 57369
rect 418 57313 486 57369
rect 542 57313 610 57369
rect 666 57313 734 57369
rect 790 57313 858 57369
rect 914 57313 982 57369
rect 1038 57313 1106 57369
rect 1162 57313 1230 57369
rect 1286 57313 1354 57369
rect 1410 57313 1478 57369
rect 1534 57313 1602 57369
rect 1658 57313 1726 57369
rect 1782 57313 1850 57369
rect 1906 57313 1916 57369
rect 104 57303 1916 57313
rect 104 56889 1916 56899
rect 104 56833 114 56889
rect 170 56833 238 56889
rect 294 56833 362 56889
rect 418 56833 486 56889
rect 542 56833 610 56889
rect 666 56833 734 56889
rect 790 56833 858 56889
rect 914 56833 982 56889
rect 1038 56833 1106 56889
rect 1162 56833 1230 56889
rect 1286 56833 1354 56889
rect 1410 56833 1478 56889
rect 1534 56833 1602 56889
rect 1658 56833 1726 56889
rect 1782 56833 1850 56889
rect 1906 56833 1916 56889
rect 104 56765 1916 56833
rect 104 56709 114 56765
rect 170 56709 238 56765
rect 294 56709 362 56765
rect 418 56709 486 56765
rect 542 56709 610 56765
rect 666 56709 734 56765
rect 790 56709 858 56765
rect 914 56709 982 56765
rect 1038 56709 1106 56765
rect 1162 56709 1230 56765
rect 1286 56709 1354 56765
rect 1410 56709 1478 56765
rect 1534 56709 1602 56765
rect 1658 56709 1726 56765
rect 1782 56709 1850 56765
rect 1906 56709 1916 56765
rect 104 56641 1916 56709
rect 104 56585 114 56641
rect 170 56585 238 56641
rect 294 56585 362 56641
rect 418 56585 486 56641
rect 542 56585 610 56641
rect 666 56585 734 56641
rect 790 56585 858 56641
rect 914 56585 982 56641
rect 1038 56585 1106 56641
rect 1162 56585 1230 56641
rect 1286 56585 1354 56641
rect 1410 56585 1478 56641
rect 1534 56585 1602 56641
rect 1658 56585 1726 56641
rect 1782 56585 1850 56641
rect 1906 56585 1916 56641
rect 104 56517 1916 56585
rect 104 56461 114 56517
rect 170 56461 238 56517
rect 294 56461 362 56517
rect 418 56461 486 56517
rect 542 56461 610 56517
rect 666 56461 734 56517
rect 790 56461 858 56517
rect 914 56461 982 56517
rect 1038 56461 1106 56517
rect 1162 56461 1230 56517
rect 1286 56461 1354 56517
rect 1410 56461 1478 56517
rect 1534 56461 1602 56517
rect 1658 56461 1726 56517
rect 1782 56461 1850 56517
rect 1906 56461 1916 56517
rect 104 56393 1916 56461
rect 104 56337 114 56393
rect 170 56337 238 56393
rect 294 56337 362 56393
rect 418 56337 486 56393
rect 542 56337 610 56393
rect 666 56337 734 56393
rect 790 56337 858 56393
rect 914 56337 982 56393
rect 1038 56337 1106 56393
rect 1162 56337 1230 56393
rect 1286 56337 1354 56393
rect 1410 56337 1478 56393
rect 1534 56337 1602 56393
rect 1658 56337 1726 56393
rect 1782 56337 1850 56393
rect 1906 56337 1916 56393
rect 104 56269 1916 56337
rect 104 56213 114 56269
rect 170 56213 238 56269
rect 294 56213 362 56269
rect 418 56213 486 56269
rect 542 56213 610 56269
rect 666 56213 734 56269
rect 790 56213 858 56269
rect 914 56213 982 56269
rect 1038 56213 1106 56269
rect 1162 56213 1230 56269
rect 1286 56213 1354 56269
rect 1410 56213 1478 56269
rect 1534 56213 1602 56269
rect 1658 56213 1726 56269
rect 1782 56213 1850 56269
rect 1906 56213 1916 56269
rect 104 56145 1916 56213
rect 104 56089 114 56145
rect 170 56089 238 56145
rect 294 56089 362 56145
rect 418 56089 486 56145
rect 542 56089 610 56145
rect 666 56089 734 56145
rect 790 56089 858 56145
rect 914 56089 982 56145
rect 1038 56089 1106 56145
rect 1162 56089 1230 56145
rect 1286 56089 1354 56145
rect 1410 56089 1478 56145
rect 1534 56089 1602 56145
rect 1658 56089 1726 56145
rect 1782 56089 1850 56145
rect 1906 56089 1916 56145
rect 104 56021 1916 56089
rect 104 55965 114 56021
rect 170 55965 238 56021
rect 294 55965 362 56021
rect 418 55965 486 56021
rect 542 55965 610 56021
rect 666 55965 734 56021
rect 790 55965 858 56021
rect 914 55965 982 56021
rect 1038 55965 1106 56021
rect 1162 55965 1230 56021
rect 1286 55965 1354 56021
rect 1410 55965 1478 56021
rect 1534 55965 1602 56021
rect 1658 55965 1726 56021
rect 1782 55965 1850 56021
rect 1906 55965 1916 56021
rect 104 55897 1916 55965
rect 104 55841 114 55897
rect 170 55841 238 55897
rect 294 55841 362 55897
rect 418 55841 486 55897
rect 542 55841 610 55897
rect 666 55841 734 55897
rect 790 55841 858 55897
rect 914 55841 982 55897
rect 1038 55841 1106 55897
rect 1162 55841 1230 55897
rect 1286 55841 1354 55897
rect 1410 55841 1478 55897
rect 1534 55841 1602 55897
rect 1658 55841 1726 55897
rect 1782 55841 1850 55897
rect 1906 55841 1916 55897
rect 104 55773 1916 55841
rect 104 55717 114 55773
rect 170 55717 238 55773
rect 294 55717 362 55773
rect 418 55717 486 55773
rect 542 55717 610 55773
rect 666 55717 734 55773
rect 790 55717 858 55773
rect 914 55717 982 55773
rect 1038 55717 1106 55773
rect 1162 55717 1230 55773
rect 1286 55717 1354 55773
rect 1410 55717 1478 55773
rect 1534 55717 1602 55773
rect 1658 55717 1726 55773
rect 1782 55717 1850 55773
rect 1906 55717 1916 55773
rect 104 55707 1916 55717
rect 104 55280 1916 55290
rect 104 55224 114 55280
rect 170 55224 238 55280
rect 294 55224 362 55280
rect 418 55224 486 55280
rect 542 55224 610 55280
rect 666 55224 734 55280
rect 790 55224 858 55280
rect 914 55224 982 55280
rect 1038 55224 1106 55280
rect 1162 55224 1230 55280
rect 1286 55224 1354 55280
rect 1410 55224 1478 55280
rect 1534 55224 1602 55280
rect 1658 55224 1726 55280
rect 1782 55224 1850 55280
rect 1906 55224 1916 55280
rect 104 55156 1916 55224
rect 104 55100 114 55156
rect 170 55100 238 55156
rect 294 55100 362 55156
rect 418 55100 486 55156
rect 542 55100 610 55156
rect 666 55100 734 55156
rect 790 55100 858 55156
rect 914 55100 982 55156
rect 1038 55100 1106 55156
rect 1162 55100 1230 55156
rect 1286 55100 1354 55156
rect 1410 55100 1478 55156
rect 1534 55100 1602 55156
rect 1658 55100 1726 55156
rect 1782 55100 1850 55156
rect 1906 55100 1916 55156
rect 104 55032 1916 55100
rect 104 54976 114 55032
rect 170 54976 238 55032
rect 294 54976 362 55032
rect 418 54976 486 55032
rect 542 54976 610 55032
rect 666 54976 734 55032
rect 790 54976 858 55032
rect 914 54976 982 55032
rect 1038 54976 1106 55032
rect 1162 54976 1230 55032
rect 1286 54976 1354 55032
rect 1410 54976 1478 55032
rect 1534 54976 1602 55032
rect 1658 54976 1726 55032
rect 1782 54976 1850 55032
rect 1906 54976 1916 55032
rect 104 54908 1916 54976
rect 104 54852 114 54908
rect 170 54852 238 54908
rect 294 54852 362 54908
rect 418 54852 486 54908
rect 542 54852 610 54908
rect 666 54852 734 54908
rect 790 54852 858 54908
rect 914 54852 982 54908
rect 1038 54852 1106 54908
rect 1162 54852 1230 54908
rect 1286 54852 1354 54908
rect 1410 54852 1478 54908
rect 1534 54852 1602 54908
rect 1658 54852 1726 54908
rect 1782 54852 1850 54908
rect 1906 54852 1916 54908
rect 104 54784 1916 54852
rect 104 54728 114 54784
rect 170 54728 238 54784
rect 294 54728 362 54784
rect 418 54728 486 54784
rect 542 54728 610 54784
rect 666 54728 734 54784
rect 790 54728 858 54784
rect 914 54728 982 54784
rect 1038 54728 1106 54784
rect 1162 54728 1230 54784
rect 1286 54728 1354 54784
rect 1410 54728 1478 54784
rect 1534 54728 1602 54784
rect 1658 54728 1726 54784
rect 1782 54728 1850 54784
rect 1906 54728 1916 54784
rect 104 54660 1916 54728
rect 104 54604 114 54660
rect 170 54604 238 54660
rect 294 54604 362 54660
rect 418 54604 486 54660
rect 542 54604 610 54660
rect 666 54604 734 54660
rect 790 54604 858 54660
rect 914 54604 982 54660
rect 1038 54604 1106 54660
rect 1162 54604 1230 54660
rect 1286 54604 1354 54660
rect 1410 54604 1478 54660
rect 1534 54604 1602 54660
rect 1658 54604 1726 54660
rect 1782 54604 1850 54660
rect 1906 54604 1916 54660
rect 104 54536 1916 54604
rect 104 54480 114 54536
rect 170 54480 238 54536
rect 294 54480 362 54536
rect 418 54480 486 54536
rect 542 54480 610 54536
rect 666 54480 734 54536
rect 790 54480 858 54536
rect 914 54480 982 54536
rect 1038 54480 1106 54536
rect 1162 54480 1230 54536
rect 1286 54480 1354 54536
rect 1410 54480 1478 54536
rect 1534 54480 1602 54536
rect 1658 54480 1726 54536
rect 1782 54480 1850 54536
rect 1906 54480 1916 54536
rect 104 54412 1916 54480
rect 104 54356 114 54412
rect 170 54356 238 54412
rect 294 54356 362 54412
rect 418 54356 486 54412
rect 542 54356 610 54412
rect 666 54356 734 54412
rect 790 54356 858 54412
rect 914 54356 982 54412
rect 1038 54356 1106 54412
rect 1162 54356 1230 54412
rect 1286 54356 1354 54412
rect 1410 54356 1478 54412
rect 1534 54356 1602 54412
rect 1658 54356 1726 54412
rect 1782 54356 1850 54412
rect 1906 54356 1916 54412
rect 104 54288 1916 54356
rect 104 54232 114 54288
rect 170 54232 238 54288
rect 294 54232 362 54288
rect 418 54232 486 54288
rect 542 54232 610 54288
rect 666 54232 734 54288
rect 790 54232 858 54288
rect 914 54232 982 54288
rect 1038 54232 1106 54288
rect 1162 54232 1230 54288
rect 1286 54232 1354 54288
rect 1410 54232 1478 54288
rect 1534 54232 1602 54288
rect 1658 54232 1726 54288
rect 1782 54232 1850 54288
rect 1906 54232 1916 54288
rect 104 54164 1916 54232
rect 104 54108 114 54164
rect 170 54108 238 54164
rect 294 54108 362 54164
rect 418 54108 486 54164
rect 542 54108 610 54164
rect 666 54108 734 54164
rect 790 54108 858 54164
rect 914 54108 982 54164
rect 1038 54108 1106 54164
rect 1162 54108 1230 54164
rect 1286 54108 1354 54164
rect 1410 54108 1478 54164
rect 1534 54108 1602 54164
rect 1658 54108 1726 54164
rect 1782 54108 1850 54164
rect 1906 54108 1916 54164
rect 104 54098 1916 54108
rect 104 53707 1916 53717
rect 104 53651 114 53707
rect 170 53651 238 53707
rect 294 53651 362 53707
rect 418 53651 486 53707
rect 542 53651 610 53707
rect 666 53651 734 53707
rect 790 53651 858 53707
rect 914 53651 982 53707
rect 1038 53651 1106 53707
rect 1162 53651 1230 53707
rect 1286 53651 1354 53707
rect 1410 53651 1478 53707
rect 1534 53651 1602 53707
rect 1658 53651 1726 53707
rect 1782 53651 1850 53707
rect 1906 53651 1916 53707
rect 104 53583 1916 53651
rect 104 53527 114 53583
rect 170 53527 238 53583
rect 294 53527 362 53583
rect 418 53527 486 53583
rect 542 53527 610 53583
rect 666 53527 734 53583
rect 790 53527 858 53583
rect 914 53527 982 53583
rect 1038 53527 1106 53583
rect 1162 53527 1230 53583
rect 1286 53527 1354 53583
rect 1410 53527 1478 53583
rect 1534 53527 1602 53583
rect 1658 53527 1726 53583
rect 1782 53527 1850 53583
rect 1906 53527 1916 53583
rect 104 53459 1916 53527
rect 104 53403 114 53459
rect 170 53403 238 53459
rect 294 53403 362 53459
rect 418 53403 486 53459
rect 542 53403 610 53459
rect 666 53403 734 53459
rect 790 53403 858 53459
rect 914 53403 982 53459
rect 1038 53403 1106 53459
rect 1162 53403 1230 53459
rect 1286 53403 1354 53459
rect 1410 53403 1478 53459
rect 1534 53403 1602 53459
rect 1658 53403 1726 53459
rect 1782 53403 1850 53459
rect 1906 53403 1916 53459
rect 104 53335 1916 53403
rect 104 53279 114 53335
rect 170 53279 238 53335
rect 294 53279 362 53335
rect 418 53279 486 53335
rect 542 53279 610 53335
rect 666 53279 734 53335
rect 790 53279 858 53335
rect 914 53279 982 53335
rect 1038 53279 1106 53335
rect 1162 53279 1230 53335
rect 1286 53279 1354 53335
rect 1410 53279 1478 53335
rect 1534 53279 1602 53335
rect 1658 53279 1726 53335
rect 1782 53279 1850 53335
rect 1906 53279 1916 53335
rect 104 53211 1916 53279
rect 104 53155 114 53211
rect 170 53155 238 53211
rect 294 53155 362 53211
rect 418 53155 486 53211
rect 542 53155 610 53211
rect 666 53155 734 53211
rect 790 53155 858 53211
rect 914 53155 982 53211
rect 1038 53155 1106 53211
rect 1162 53155 1230 53211
rect 1286 53155 1354 53211
rect 1410 53155 1478 53211
rect 1534 53155 1602 53211
rect 1658 53155 1726 53211
rect 1782 53155 1850 53211
rect 1906 53155 1916 53211
rect 104 53087 1916 53155
rect 104 53031 114 53087
rect 170 53031 238 53087
rect 294 53031 362 53087
rect 418 53031 486 53087
rect 542 53031 610 53087
rect 666 53031 734 53087
rect 790 53031 858 53087
rect 914 53031 982 53087
rect 1038 53031 1106 53087
rect 1162 53031 1230 53087
rect 1286 53031 1354 53087
rect 1410 53031 1478 53087
rect 1534 53031 1602 53087
rect 1658 53031 1726 53087
rect 1782 53031 1850 53087
rect 1906 53031 1916 53087
rect 104 52963 1916 53031
rect 104 52907 114 52963
rect 170 52907 238 52963
rect 294 52907 362 52963
rect 418 52907 486 52963
rect 542 52907 610 52963
rect 666 52907 734 52963
rect 790 52907 858 52963
rect 914 52907 982 52963
rect 1038 52907 1106 52963
rect 1162 52907 1230 52963
rect 1286 52907 1354 52963
rect 1410 52907 1478 52963
rect 1534 52907 1602 52963
rect 1658 52907 1726 52963
rect 1782 52907 1850 52963
rect 1906 52907 1916 52963
rect 104 52839 1916 52907
rect 104 52783 114 52839
rect 170 52783 238 52839
rect 294 52783 362 52839
rect 418 52783 486 52839
rect 542 52783 610 52839
rect 666 52783 734 52839
rect 790 52783 858 52839
rect 914 52783 982 52839
rect 1038 52783 1106 52839
rect 1162 52783 1230 52839
rect 1286 52783 1354 52839
rect 1410 52783 1478 52839
rect 1534 52783 1602 52839
rect 1658 52783 1726 52839
rect 1782 52783 1850 52839
rect 1906 52783 1916 52839
rect 104 52715 1916 52783
rect 104 52659 114 52715
rect 170 52659 238 52715
rect 294 52659 362 52715
rect 418 52659 486 52715
rect 542 52659 610 52715
rect 666 52659 734 52715
rect 790 52659 858 52715
rect 914 52659 982 52715
rect 1038 52659 1106 52715
rect 1162 52659 1230 52715
rect 1286 52659 1354 52715
rect 1410 52659 1478 52715
rect 1534 52659 1602 52715
rect 1658 52659 1726 52715
rect 1782 52659 1850 52715
rect 1906 52659 1916 52715
rect 104 52591 1916 52659
rect 104 52535 114 52591
rect 170 52535 238 52591
rect 294 52535 362 52591
rect 418 52535 486 52591
rect 542 52535 610 52591
rect 666 52535 734 52591
rect 790 52535 858 52591
rect 914 52535 982 52591
rect 1038 52535 1106 52591
rect 1162 52535 1230 52591
rect 1286 52535 1354 52591
rect 1410 52535 1478 52591
rect 1534 52535 1602 52591
rect 1658 52535 1726 52591
rect 1782 52535 1850 52591
rect 1906 52535 1916 52591
rect 104 52525 1916 52535
rect 104 52100 1916 52110
rect 104 52044 114 52100
rect 170 52044 238 52100
rect 294 52044 362 52100
rect 418 52044 486 52100
rect 542 52044 610 52100
rect 666 52044 734 52100
rect 790 52044 858 52100
rect 914 52044 982 52100
rect 1038 52044 1106 52100
rect 1162 52044 1230 52100
rect 1286 52044 1354 52100
rect 1410 52044 1478 52100
rect 1534 52044 1602 52100
rect 1658 52044 1726 52100
rect 1782 52044 1850 52100
rect 1906 52044 1916 52100
rect 104 51976 1916 52044
rect 104 51920 114 51976
rect 170 51920 238 51976
rect 294 51920 362 51976
rect 418 51920 486 51976
rect 542 51920 610 51976
rect 666 51920 734 51976
rect 790 51920 858 51976
rect 914 51920 982 51976
rect 1038 51920 1106 51976
rect 1162 51920 1230 51976
rect 1286 51920 1354 51976
rect 1410 51920 1478 51976
rect 1534 51920 1602 51976
rect 1658 51920 1726 51976
rect 1782 51920 1850 51976
rect 1906 51920 1916 51976
rect 104 51852 1916 51920
rect 104 51796 114 51852
rect 170 51796 238 51852
rect 294 51796 362 51852
rect 418 51796 486 51852
rect 542 51796 610 51852
rect 666 51796 734 51852
rect 790 51796 858 51852
rect 914 51796 982 51852
rect 1038 51796 1106 51852
rect 1162 51796 1230 51852
rect 1286 51796 1354 51852
rect 1410 51796 1478 51852
rect 1534 51796 1602 51852
rect 1658 51796 1726 51852
rect 1782 51796 1850 51852
rect 1906 51796 1916 51852
rect 104 51728 1916 51796
rect 104 51672 114 51728
rect 170 51672 238 51728
rect 294 51672 362 51728
rect 418 51672 486 51728
rect 542 51672 610 51728
rect 666 51672 734 51728
rect 790 51672 858 51728
rect 914 51672 982 51728
rect 1038 51672 1106 51728
rect 1162 51672 1230 51728
rect 1286 51672 1354 51728
rect 1410 51672 1478 51728
rect 1534 51672 1602 51728
rect 1658 51672 1726 51728
rect 1782 51672 1850 51728
rect 1906 51672 1916 51728
rect 104 51604 1916 51672
rect 104 51548 114 51604
rect 170 51548 238 51604
rect 294 51548 362 51604
rect 418 51548 486 51604
rect 542 51548 610 51604
rect 666 51548 734 51604
rect 790 51548 858 51604
rect 914 51548 982 51604
rect 1038 51548 1106 51604
rect 1162 51548 1230 51604
rect 1286 51548 1354 51604
rect 1410 51548 1478 51604
rect 1534 51548 1602 51604
rect 1658 51548 1726 51604
rect 1782 51548 1850 51604
rect 1906 51548 1916 51604
rect 104 51480 1916 51548
rect 104 51424 114 51480
rect 170 51424 238 51480
rect 294 51424 362 51480
rect 418 51424 486 51480
rect 542 51424 610 51480
rect 666 51424 734 51480
rect 790 51424 858 51480
rect 914 51424 982 51480
rect 1038 51424 1106 51480
rect 1162 51424 1230 51480
rect 1286 51424 1354 51480
rect 1410 51424 1478 51480
rect 1534 51424 1602 51480
rect 1658 51424 1726 51480
rect 1782 51424 1850 51480
rect 1906 51424 1916 51480
rect 104 51356 1916 51424
rect 104 51300 114 51356
rect 170 51300 238 51356
rect 294 51300 362 51356
rect 418 51300 486 51356
rect 542 51300 610 51356
rect 666 51300 734 51356
rect 790 51300 858 51356
rect 914 51300 982 51356
rect 1038 51300 1106 51356
rect 1162 51300 1230 51356
rect 1286 51300 1354 51356
rect 1410 51300 1478 51356
rect 1534 51300 1602 51356
rect 1658 51300 1726 51356
rect 1782 51300 1850 51356
rect 1906 51300 1916 51356
rect 104 51232 1916 51300
rect 104 51176 114 51232
rect 170 51176 238 51232
rect 294 51176 362 51232
rect 418 51176 486 51232
rect 542 51176 610 51232
rect 666 51176 734 51232
rect 790 51176 858 51232
rect 914 51176 982 51232
rect 1038 51176 1106 51232
rect 1162 51176 1230 51232
rect 1286 51176 1354 51232
rect 1410 51176 1478 51232
rect 1534 51176 1602 51232
rect 1658 51176 1726 51232
rect 1782 51176 1850 51232
rect 1906 51176 1916 51232
rect 104 51108 1916 51176
rect 104 51052 114 51108
rect 170 51052 238 51108
rect 294 51052 362 51108
rect 418 51052 486 51108
rect 542 51052 610 51108
rect 666 51052 734 51108
rect 790 51052 858 51108
rect 914 51052 982 51108
rect 1038 51052 1106 51108
rect 1162 51052 1230 51108
rect 1286 51052 1354 51108
rect 1410 51052 1478 51108
rect 1534 51052 1602 51108
rect 1658 51052 1726 51108
rect 1782 51052 1850 51108
rect 1906 51052 1916 51108
rect 104 50984 1916 51052
rect 104 50928 114 50984
rect 170 50928 238 50984
rect 294 50928 362 50984
rect 418 50928 486 50984
rect 542 50928 610 50984
rect 666 50928 734 50984
rect 790 50928 858 50984
rect 914 50928 982 50984
rect 1038 50928 1106 50984
rect 1162 50928 1230 50984
rect 1286 50928 1354 50984
rect 1410 50928 1478 50984
rect 1534 50928 1602 50984
rect 1658 50928 1726 50984
rect 1782 50928 1850 50984
rect 1906 50928 1916 50984
rect 104 50918 1916 50928
rect 104 50480 1916 50490
rect 104 50424 114 50480
rect 170 50424 238 50480
rect 294 50424 362 50480
rect 418 50424 486 50480
rect 542 50424 610 50480
rect 666 50424 734 50480
rect 790 50424 858 50480
rect 914 50424 982 50480
rect 1038 50424 1106 50480
rect 1162 50424 1230 50480
rect 1286 50424 1354 50480
rect 1410 50424 1478 50480
rect 1534 50424 1602 50480
rect 1658 50424 1726 50480
rect 1782 50424 1850 50480
rect 1906 50424 1916 50480
rect 104 50356 1916 50424
rect 104 50300 114 50356
rect 170 50300 238 50356
rect 294 50300 362 50356
rect 418 50300 486 50356
rect 542 50300 610 50356
rect 666 50300 734 50356
rect 790 50300 858 50356
rect 914 50300 982 50356
rect 1038 50300 1106 50356
rect 1162 50300 1230 50356
rect 1286 50300 1354 50356
rect 1410 50300 1478 50356
rect 1534 50300 1602 50356
rect 1658 50300 1726 50356
rect 1782 50300 1850 50356
rect 1906 50300 1916 50356
rect 104 50232 1916 50300
rect 104 50176 114 50232
rect 170 50176 238 50232
rect 294 50176 362 50232
rect 418 50176 486 50232
rect 542 50176 610 50232
rect 666 50176 734 50232
rect 790 50176 858 50232
rect 914 50176 982 50232
rect 1038 50176 1106 50232
rect 1162 50176 1230 50232
rect 1286 50176 1354 50232
rect 1410 50176 1478 50232
rect 1534 50176 1602 50232
rect 1658 50176 1726 50232
rect 1782 50176 1850 50232
rect 1906 50176 1916 50232
rect 104 50108 1916 50176
rect 104 50052 114 50108
rect 170 50052 238 50108
rect 294 50052 362 50108
rect 418 50052 486 50108
rect 542 50052 610 50108
rect 666 50052 734 50108
rect 790 50052 858 50108
rect 914 50052 982 50108
rect 1038 50052 1106 50108
rect 1162 50052 1230 50108
rect 1286 50052 1354 50108
rect 1410 50052 1478 50108
rect 1534 50052 1602 50108
rect 1658 50052 1726 50108
rect 1782 50052 1850 50108
rect 1906 50052 1916 50108
rect 104 49984 1916 50052
rect 104 49928 114 49984
rect 170 49928 238 49984
rect 294 49928 362 49984
rect 418 49928 486 49984
rect 542 49928 610 49984
rect 666 49928 734 49984
rect 790 49928 858 49984
rect 914 49928 982 49984
rect 1038 49928 1106 49984
rect 1162 49928 1230 49984
rect 1286 49928 1354 49984
rect 1410 49928 1478 49984
rect 1534 49928 1602 49984
rect 1658 49928 1726 49984
rect 1782 49928 1850 49984
rect 1906 49928 1916 49984
rect 104 49860 1916 49928
rect 104 49804 114 49860
rect 170 49804 238 49860
rect 294 49804 362 49860
rect 418 49804 486 49860
rect 542 49804 610 49860
rect 666 49804 734 49860
rect 790 49804 858 49860
rect 914 49804 982 49860
rect 1038 49804 1106 49860
rect 1162 49804 1230 49860
rect 1286 49804 1354 49860
rect 1410 49804 1478 49860
rect 1534 49804 1602 49860
rect 1658 49804 1726 49860
rect 1782 49804 1850 49860
rect 1906 49804 1916 49860
rect 104 49736 1916 49804
rect 104 49680 114 49736
rect 170 49680 238 49736
rect 294 49680 362 49736
rect 418 49680 486 49736
rect 542 49680 610 49736
rect 666 49680 734 49736
rect 790 49680 858 49736
rect 914 49680 982 49736
rect 1038 49680 1106 49736
rect 1162 49680 1230 49736
rect 1286 49680 1354 49736
rect 1410 49680 1478 49736
rect 1534 49680 1602 49736
rect 1658 49680 1726 49736
rect 1782 49680 1850 49736
rect 1906 49680 1916 49736
rect 104 49612 1916 49680
rect 104 49556 114 49612
rect 170 49556 238 49612
rect 294 49556 362 49612
rect 418 49556 486 49612
rect 542 49556 610 49612
rect 666 49556 734 49612
rect 790 49556 858 49612
rect 914 49556 982 49612
rect 1038 49556 1106 49612
rect 1162 49556 1230 49612
rect 1286 49556 1354 49612
rect 1410 49556 1478 49612
rect 1534 49556 1602 49612
rect 1658 49556 1726 49612
rect 1782 49556 1850 49612
rect 1906 49556 1916 49612
rect 104 49488 1916 49556
rect 104 49432 114 49488
rect 170 49432 238 49488
rect 294 49432 362 49488
rect 418 49432 486 49488
rect 542 49432 610 49488
rect 666 49432 734 49488
rect 790 49432 858 49488
rect 914 49432 982 49488
rect 1038 49432 1106 49488
rect 1162 49432 1230 49488
rect 1286 49432 1354 49488
rect 1410 49432 1478 49488
rect 1534 49432 1602 49488
rect 1658 49432 1726 49488
rect 1782 49432 1850 49488
rect 1906 49432 1916 49488
rect 104 49364 1916 49432
rect 104 49308 114 49364
rect 170 49308 238 49364
rect 294 49308 362 49364
rect 418 49308 486 49364
rect 542 49308 610 49364
rect 666 49308 734 49364
rect 790 49308 858 49364
rect 914 49308 982 49364
rect 1038 49308 1106 49364
rect 1162 49308 1230 49364
rect 1286 49308 1354 49364
rect 1410 49308 1478 49364
rect 1534 49308 1602 49364
rect 1658 49308 1726 49364
rect 1782 49308 1850 49364
rect 1906 49308 1916 49364
rect 104 49298 1916 49308
rect 104 48841 1916 48851
rect 104 48785 114 48841
rect 170 48785 238 48841
rect 294 48785 362 48841
rect 418 48785 486 48841
rect 542 48785 610 48841
rect 666 48785 734 48841
rect 790 48785 858 48841
rect 914 48785 982 48841
rect 1038 48785 1106 48841
rect 1162 48785 1230 48841
rect 1286 48785 1354 48841
rect 1410 48785 1478 48841
rect 1534 48785 1602 48841
rect 1658 48785 1726 48841
rect 1782 48785 1850 48841
rect 1906 48785 1916 48841
rect 104 48717 1916 48785
rect 104 48661 114 48717
rect 170 48661 238 48717
rect 294 48661 362 48717
rect 418 48661 486 48717
rect 542 48661 610 48717
rect 666 48661 734 48717
rect 790 48661 858 48717
rect 914 48661 982 48717
rect 1038 48661 1106 48717
rect 1162 48661 1230 48717
rect 1286 48661 1354 48717
rect 1410 48661 1478 48717
rect 1534 48661 1602 48717
rect 1658 48661 1726 48717
rect 1782 48661 1850 48717
rect 1906 48661 1916 48717
rect 104 48593 1916 48661
rect 104 48537 114 48593
rect 170 48537 238 48593
rect 294 48537 362 48593
rect 418 48537 486 48593
rect 542 48537 610 48593
rect 666 48537 734 48593
rect 790 48537 858 48593
rect 914 48537 982 48593
rect 1038 48537 1106 48593
rect 1162 48537 1230 48593
rect 1286 48537 1354 48593
rect 1410 48537 1478 48593
rect 1534 48537 1602 48593
rect 1658 48537 1726 48593
rect 1782 48537 1850 48593
rect 1906 48537 1916 48593
rect 104 48469 1916 48537
rect 104 48413 114 48469
rect 170 48413 238 48469
rect 294 48413 362 48469
rect 418 48413 486 48469
rect 542 48413 610 48469
rect 666 48413 734 48469
rect 790 48413 858 48469
rect 914 48413 982 48469
rect 1038 48413 1106 48469
rect 1162 48413 1230 48469
rect 1286 48413 1354 48469
rect 1410 48413 1478 48469
rect 1534 48413 1602 48469
rect 1658 48413 1726 48469
rect 1782 48413 1850 48469
rect 1906 48413 1916 48469
rect 104 48345 1916 48413
rect 104 48289 114 48345
rect 170 48289 238 48345
rect 294 48289 362 48345
rect 418 48289 486 48345
rect 542 48289 610 48345
rect 666 48289 734 48345
rect 790 48289 858 48345
rect 914 48289 982 48345
rect 1038 48289 1106 48345
rect 1162 48289 1230 48345
rect 1286 48289 1354 48345
rect 1410 48289 1478 48345
rect 1534 48289 1602 48345
rect 1658 48289 1726 48345
rect 1782 48289 1850 48345
rect 1906 48289 1916 48345
rect 104 48221 1916 48289
rect 104 48165 114 48221
rect 170 48165 238 48221
rect 294 48165 362 48221
rect 418 48165 486 48221
rect 542 48165 610 48221
rect 666 48165 734 48221
rect 790 48165 858 48221
rect 914 48165 982 48221
rect 1038 48165 1106 48221
rect 1162 48165 1230 48221
rect 1286 48165 1354 48221
rect 1410 48165 1478 48221
rect 1534 48165 1602 48221
rect 1658 48165 1726 48221
rect 1782 48165 1850 48221
rect 1906 48165 1916 48221
rect 104 48097 1916 48165
rect 104 48041 114 48097
rect 170 48041 238 48097
rect 294 48041 362 48097
rect 418 48041 486 48097
rect 542 48041 610 48097
rect 666 48041 734 48097
rect 790 48041 858 48097
rect 914 48041 982 48097
rect 1038 48041 1106 48097
rect 1162 48041 1230 48097
rect 1286 48041 1354 48097
rect 1410 48041 1478 48097
rect 1534 48041 1602 48097
rect 1658 48041 1726 48097
rect 1782 48041 1850 48097
rect 1906 48041 1916 48097
rect 104 47973 1916 48041
rect 104 47917 114 47973
rect 170 47917 238 47973
rect 294 47917 362 47973
rect 418 47917 486 47973
rect 542 47917 610 47973
rect 666 47917 734 47973
rect 790 47917 858 47973
rect 914 47917 982 47973
rect 1038 47917 1106 47973
rect 1162 47917 1230 47973
rect 1286 47917 1354 47973
rect 1410 47917 1478 47973
rect 1534 47917 1602 47973
rect 1658 47917 1726 47973
rect 1782 47917 1850 47973
rect 1906 47917 1916 47973
rect 104 47849 1916 47917
rect 104 47793 114 47849
rect 170 47793 238 47849
rect 294 47793 362 47849
rect 418 47793 486 47849
rect 542 47793 610 47849
rect 666 47793 734 47849
rect 790 47793 858 47849
rect 914 47793 982 47849
rect 1038 47793 1106 47849
rect 1162 47793 1230 47849
rect 1286 47793 1354 47849
rect 1410 47793 1478 47849
rect 1534 47793 1602 47849
rect 1658 47793 1726 47849
rect 1782 47793 1850 47849
rect 1906 47793 1916 47849
rect 104 47725 1916 47793
rect 104 47669 114 47725
rect 170 47669 238 47725
rect 294 47669 362 47725
rect 418 47669 486 47725
rect 542 47669 610 47725
rect 666 47669 734 47725
rect 790 47669 858 47725
rect 914 47669 982 47725
rect 1038 47669 1106 47725
rect 1162 47669 1230 47725
rect 1286 47669 1354 47725
rect 1410 47669 1478 47725
rect 1534 47669 1602 47725
rect 1658 47669 1726 47725
rect 1782 47669 1850 47725
rect 1906 47669 1916 47725
rect 104 47601 1916 47669
rect 104 47545 114 47601
rect 170 47545 238 47601
rect 294 47545 362 47601
rect 418 47545 486 47601
rect 542 47545 610 47601
rect 666 47545 734 47601
rect 790 47545 858 47601
rect 914 47545 982 47601
rect 1038 47545 1106 47601
rect 1162 47545 1230 47601
rect 1286 47545 1354 47601
rect 1410 47545 1478 47601
rect 1534 47545 1602 47601
rect 1658 47545 1726 47601
rect 1782 47545 1850 47601
rect 1906 47545 1916 47601
rect 104 47477 1916 47545
rect 104 47421 114 47477
rect 170 47421 238 47477
rect 294 47421 362 47477
rect 418 47421 486 47477
rect 542 47421 610 47477
rect 666 47421 734 47477
rect 790 47421 858 47477
rect 914 47421 982 47477
rect 1038 47421 1106 47477
rect 1162 47421 1230 47477
rect 1286 47421 1354 47477
rect 1410 47421 1478 47477
rect 1534 47421 1602 47477
rect 1658 47421 1726 47477
rect 1782 47421 1850 47477
rect 1906 47421 1916 47477
rect 104 47353 1916 47421
rect 104 47297 114 47353
rect 170 47297 238 47353
rect 294 47297 362 47353
rect 418 47297 486 47353
rect 542 47297 610 47353
rect 666 47297 734 47353
rect 790 47297 858 47353
rect 914 47297 982 47353
rect 1038 47297 1106 47353
rect 1162 47297 1230 47353
rect 1286 47297 1354 47353
rect 1410 47297 1478 47353
rect 1534 47297 1602 47353
rect 1658 47297 1726 47353
rect 1782 47297 1850 47353
rect 1906 47297 1916 47353
rect 104 47229 1916 47297
rect 104 47173 114 47229
rect 170 47173 238 47229
rect 294 47173 362 47229
rect 418 47173 486 47229
rect 542 47173 610 47229
rect 666 47173 734 47229
rect 790 47173 858 47229
rect 914 47173 982 47229
rect 1038 47173 1106 47229
rect 1162 47173 1230 47229
rect 1286 47173 1354 47229
rect 1410 47173 1478 47229
rect 1534 47173 1602 47229
rect 1658 47173 1726 47229
rect 1782 47173 1850 47229
rect 1906 47173 1916 47229
rect 104 47105 1916 47173
rect 104 47049 114 47105
rect 170 47049 238 47105
rect 294 47049 362 47105
rect 418 47049 486 47105
rect 542 47049 610 47105
rect 666 47049 734 47105
rect 790 47049 858 47105
rect 914 47049 982 47105
rect 1038 47049 1106 47105
rect 1162 47049 1230 47105
rect 1286 47049 1354 47105
rect 1410 47049 1478 47105
rect 1534 47049 1602 47105
rect 1658 47049 1726 47105
rect 1782 47049 1850 47105
rect 1906 47049 1916 47105
rect 104 46981 1916 47049
rect 104 46925 114 46981
rect 170 46925 238 46981
rect 294 46925 362 46981
rect 418 46925 486 46981
rect 542 46925 610 46981
rect 666 46925 734 46981
rect 790 46925 858 46981
rect 914 46925 982 46981
rect 1038 46925 1106 46981
rect 1162 46925 1230 46981
rect 1286 46925 1354 46981
rect 1410 46925 1478 46981
rect 1534 46925 1602 46981
rect 1658 46925 1726 46981
rect 1782 46925 1850 46981
rect 1906 46925 1916 46981
rect 104 46857 1916 46925
rect 104 46801 114 46857
rect 170 46801 238 46857
rect 294 46801 362 46857
rect 418 46801 486 46857
rect 542 46801 610 46857
rect 666 46801 734 46857
rect 790 46801 858 46857
rect 914 46801 982 46857
rect 1038 46801 1106 46857
rect 1162 46801 1230 46857
rect 1286 46801 1354 46857
rect 1410 46801 1478 46857
rect 1534 46801 1602 46857
rect 1658 46801 1726 46857
rect 1782 46801 1850 46857
rect 1906 46801 1916 46857
rect 104 46733 1916 46801
rect 104 46677 114 46733
rect 170 46677 238 46733
rect 294 46677 362 46733
rect 418 46677 486 46733
rect 542 46677 610 46733
rect 666 46677 734 46733
rect 790 46677 858 46733
rect 914 46677 982 46733
rect 1038 46677 1106 46733
rect 1162 46677 1230 46733
rect 1286 46677 1354 46733
rect 1410 46677 1478 46733
rect 1534 46677 1602 46733
rect 1658 46677 1726 46733
rect 1782 46677 1850 46733
rect 1906 46677 1916 46733
rect 104 46609 1916 46677
rect 104 46553 114 46609
rect 170 46553 238 46609
rect 294 46553 362 46609
rect 418 46553 486 46609
rect 542 46553 610 46609
rect 666 46553 734 46609
rect 790 46553 858 46609
rect 914 46553 982 46609
rect 1038 46553 1106 46609
rect 1162 46553 1230 46609
rect 1286 46553 1354 46609
rect 1410 46553 1478 46609
rect 1534 46553 1602 46609
rect 1658 46553 1726 46609
rect 1782 46553 1850 46609
rect 1906 46553 1916 46609
rect 104 46485 1916 46553
rect 104 46429 114 46485
rect 170 46429 238 46485
rect 294 46429 362 46485
rect 418 46429 486 46485
rect 542 46429 610 46485
rect 666 46429 734 46485
rect 790 46429 858 46485
rect 914 46429 982 46485
rect 1038 46429 1106 46485
rect 1162 46429 1230 46485
rect 1286 46429 1354 46485
rect 1410 46429 1478 46485
rect 1534 46429 1602 46485
rect 1658 46429 1726 46485
rect 1782 46429 1850 46485
rect 1906 46429 1916 46485
rect 104 46361 1916 46429
rect 104 46305 114 46361
rect 170 46305 238 46361
rect 294 46305 362 46361
rect 418 46305 486 46361
rect 542 46305 610 46361
rect 666 46305 734 46361
rect 790 46305 858 46361
rect 914 46305 982 46361
rect 1038 46305 1106 46361
rect 1162 46305 1230 46361
rect 1286 46305 1354 46361
rect 1410 46305 1478 46361
rect 1534 46305 1602 46361
rect 1658 46305 1726 46361
rect 1782 46305 1850 46361
rect 1906 46305 1916 46361
rect 104 46237 1916 46305
rect 104 46181 114 46237
rect 170 46181 238 46237
rect 294 46181 362 46237
rect 418 46181 486 46237
rect 542 46181 610 46237
rect 666 46181 734 46237
rect 790 46181 858 46237
rect 914 46181 982 46237
rect 1038 46181 1106 46237
rect 1162 46181 1230 46237
rect 1286 46181 1354 46237
rect 1410 46181 1478 46237
rect 1534 46181 1602 46237
rect 1658 46181 1726 46237
rect 1782 46181 1850 46237
rect 1906 46181 1916 46237
rect 104 46171 1916 46181
rect 104 45652 1916 45662
rect 104 45596 114 45652
rect 170 45596 238 45652
rect 294 45596 362 45652
rect 418 45596 486 45652
rect 542 45596 610 45652
rect 666 45596 734 45652
rect 790 45596 858 45652
rect 914 45596 982 45652
rect 1038 45596 1106 45652
rect 1162 45596 1230 45652
rect 1286 45596 1354 45652
rect 1410 45596 1478 45652
rect 1534 45596 1602 45652
rect 1658 45596 1726 45652
rect 1782 45596 1850 45652
rect 1906 45596 1916 45652
rect 104 45528 1916 45596
rect 104 45472 114 45528
rect 170 45472 238 45528
rect 294 45472 362 45528
rect 418 45472 486 45528
rect 542 45472 610 45528
rect 666 45472 734 45528
rect 790 45472 858 45528
rect 914 45472 982 45528
rect 1038 45472 1106 45528
rect 1162 45472 1230 45528
rect 1286 45472 1354 45528
rect 1410 45472 1478 45528
rect 1534 45472 1602 45528
rect 1658 45472 1726 45528
rect 1782 45472 1850 45528
rect 1906 45472 1916 45528
rect 104 45404 1916 45472
rect 104 45348 114 45404
rect 170 45348 238 45404
rect 294 45348 362 45404
rect 418 45348 486 45404
rect 542 45348 610 45404
rect 666 45348 734 45404
rect 790 45348 858 45404
rect 914 45348 982 45404
rect 1038 45348 1106 45404
rect 1162 45348 1230 45404
rect 1286 45348 1354 45404
rect 1410 45348 1478 45404
rect 1534 45348 1602 45404
rect 1658 45348 1726 45404
rect 1782 45348 1850 45404
rect 1906 45348 1916 45404
rect 104 45280 1916 45348
rect 104 45224 114 45280
rect 170 45224 238 45280
rect 294 45224 362 45280
rect 418 45224 486 45280
rect 542 45224 610 45280
rect 666 45224 734 45280
rect 790 45224 858 45280
rect 914 45224 982 45280
rect 1038 45224 1106 45280
rect 1162 45224 1230 45280
rect 1286 45224 1354 45280
rect 1410 45224 1478 45280
rect 1534 45224 1602 45280
rect 1658 45224 1726 45280
rect 1782 45224 1850 45280
rect 1906 45224 1916 45280
rect 104 45156 1916 45224
rect 104 45100 114 45156
rect 170 45100 238 45156
rect 294 45100 362 45156
rect 418 45100 486 45156
rect 542 45100 610 45156
rect 666 45100 734 45156
rect 790 45100 858 45156
rect 914 45100 982 45156
rect 1038 45100 1106 45156
rect 1162 45100 1230 45156
rect 1286 45100 1354 45156
rect 1410 45100 1478 45156
rect 1534 45100 1602 45156
rect 1658 45100 1726 45156
rect 1782 45100 1850 45156
rect 1906 45100 1916 45156
rect 104 45032 1916 45100
rect 104 44976 114 45032
rect 170 44976 238 45032
rect 294 44976 362 45032
rect 418 44976 486 45032
rect 542 44976 610 45032
rect 666 44976 734 45032
rect 790 44976 858 45032
rect 914 44976 982 45032
rect 1038 44976 1106 45032
rect 1162 44976 1230 45032
rect 1286 44976 1354 45032
rect 1410 44976 1478 45032
rect 1534 44976 1602 45032
rect 1658 44976 1726 45032
rect 1782 44976 1850 45032
rect 1906 44976 1916 45032
rect 104 44908 1916 44976
rect 104 44852 114 44908
rect 170 44852 238 44908
rect 294 44852 362 44908
rect 418 44852 486 44908
rect 542 44852 610 44908
rect 666 44852 734 44908
rect 790 44852 858 44908
rect 914 44852 982 44908
rect 1038 44852 1106 44908
rect 1162 44852 1230 44908
rect 1286 44852 1354 44908
rect 1410 44852 1478 44908
rect 1534 44852 1602 44908
rect 1658 44852 1726 44908
rect 1782 44852 1850 44908
rect 1906 44852 1916 44908
rect 104 44784 1916 44852
rect 104 44728 114 44784
rect 170 44728 238 44784
rect 294 44728 362 44784
rect 418 44728 486 44784
rect 542 44728 610 44784
rect 666 44728 734 44784
rect 790 44728 858 44784
rect 914 44728 982 44784
rect 1038 44728 1106 44784
rect 1162 44728 1230 44784
rect 1286 44728 1354 44784
rect 1410 44728 1478 44784
rect 1534 44728 1602 44784
rect 1658 44728 1726 44784
rect 1782 44728 1850 44784
rect 1906 44728 1916 44784
rect 104 44660 1916 44728
rect 104 44604 114 44660
rect 170 44604 238 44660
rect 294 44604 362 44660
rect 418 44604 486 44660
rect 542 44604 610 44660
rect 666 44604 734 44660
rect 790 44604 858 44660
rect 914 44604 982 44660
rect 1038 44604 1106 44660
rect 1162 44604 1230 44660
rect 1286 44604 1354 44660
rect 1410 44604 1478 44660
rect 1534 44604 1602 44660
rect 1658 44604 1726 44660
rect 1782 44604 1850 44660
rect 1906 44604 1916 44660
rect 104 44536 1916 44604
rect 104 44480 114 44536
rect 170 44480 238 44536
rect 294 44480 362 44536
rect 418 44480 486 44536
rect 542 44480 610 44536
rect 666 44480 734 44536
rect 790 44480 858 44536
rect 914 44480 982 44536
rect 1038 44480 1106 44536
rect 1162 44480 1230 44536
rect 1286 44480 1354 44536
rect 1410 44480 1478 44536
rect 1534 44480 1602 44536
rect 1658 44480 1726 44536
rect 1782 44480 1850 44536
rect 1906 44480 1916 44536
rect 104 44412 1916 44480
rect 104 44356 114 44412
rect 170 44356 238 44412
rect 294 44356 362 44412
rect 418 44356 486 44412
rect 542 44356 610 44412
rect 666 44356 734 44412
rect 790 44356 858 44412
rect 914 44356 982 44412
rect 1038 44356 1106 44412
rect 1162 44356 1230 44412
rect 1286 44356 1354 44412
rect 1410 44356 1478 44412
rect 1534 44356 1602 44412
rect 1658 44356 1726 44412
rect 1782 44356 1850 44412
rect 1906 44356 1916 44412
rect 104 44288 1916 44356
rect 104 44232 114 44288
rect 170 44232 238 44288
rect 294 44232 362 44288
rect 418 44232 486 44288
rect 542 44232 610 44288
rect 666 44232 734 44288
rect 790 44232 858 44288
rect 914 44232 982 44288
rect 1038 44232 1106 44288
rect 1162 44232 1230 44288
rect 1286 44232 1354 44288
rect 1410 44232 1478 44288
rect 1534 44232 1602 44288
rect 1658 44232 1726 44288
rect 1782 44232 1850 44288
rect 1906 44232 1916 44288
rect 104 44164 1916 44232
rect 104 44108 114 44164
rect 170 44108 238 44164
rect 294 44108 362 44164
rect 418 44108 486 44164
rect 542 44108 610 44164
rect 666 44108 734 44164
rect 790 44108 858 44164
rect 914 44108 982 44164
rect 1038 44108 1106 44164
rect 1162 44108 1230 44164
rect 1286 44108 1354 44164
rect 1410 44108 1478 44164
rect 1534 44108 1602 44164
rect 1658 44108 1726 44164
rect 1782 44108 1850 44164
rect 1906 44108 1916 44164
rect 104 44040 1916 44108
rect 104 43984 114 44040
rect 170 43984 238 44040
rect 294 43984 362 44040
rect 418 43984 486 44040
rect 542 43984 610 44040
rect 666 43984 734 44040
rect 790 43984 858 44040
rect 914 43984 982 44040
rect 1038 43984 1106 44040
rect 1162 43984 1230 44040
rect 1286 43984 1354 44040
rect 1410 43984 1478 44040
rect 1534 43984 1602 44040
rect 1658 43984 1726 44040
rect 1782 43984 1850 44040
rect 1906 43984 1916 44040
rect 104 43916 1916 43984
rect 104 43860 114 43916
rect 170 43860 238 43916
rect 294 43860 362 43916
rect 418 43860 486 43916
rect 542 43860 610 43916
rect 666 43860 734 43916
rect 790 43860 858 43916
rect 914 43860 982 43916
rect 1038 43860 1106 43916
rect 1162 43860 1230 43916
rect 1286 43860 1354 43916
rect 1410 43860 1478 43916
rect 1534 43860 1602 43916
rect 1658 43860 1726 43916
rect 1782 43860 1850 43916
rect 1906 43860 1916 43916
rect 104 43792 1916 43860
rect 104 43736 114 43792
rect 170 43736 238 43792
rect 294 43736 362 43792
rect 418 43736 486 43792
rect 542 43736 610 43792
rect 666 43736 734 43792
rect 790 43736 858 43792
rect 914 43736 982 43792
rect 1038 43736 1106 43792
rect 1162 43736 1230 43792
rect 1286 43736 1354 43792
rect 1410 43736 1478 43792
rect 1534 43736 1602 43792
rect 1658 43736 1726 43792
rect 1782 43736 1850 43792
rect 1906 43736 1916 43792
rect 104 43668 1916 43736
rect 104 43612 114 43668
rect 170 43612 238 43668
rect 294 43612 362 43668
rect 418 43612 486 43668
rect 542 43612 610 43668
rect 666 43612 734 43668
rect 790 43612 858 43668
rect 914 43612 982 43668
rect 1038 43612 1106 43668
rect 1162 43612 1230 43668
rect 1286 43612 1354 43668
rect 1410 43612 1478 43668
rect 1534 43612 1602 43668
rect 1658 43612 1726 43668
rect 1782 43612 1850 43668
rect 1906 43612 1916 43668
rect 104 43544 1916 43612
rect 104 43488 114 43544
rect 170 43488 238 43544
rect 294 43488 362 43544
rect 418 43488 486 43544
rect 542 43488 610 43544
rect 666 43488 734 43544
rect 790 43488 858 43544
rect 914 43488 982 43544
rect 1038 43488 1106 43544
rect 1162 43488 1230 43544
rect 1286 43488 1354 43544
rect 1410 43488 1478 43544
rect 1534 43488 1602 43544
rect 1658 43488 1726 43544
rect 1782 43488 1850 43544
rect 1906 43488 1916 43544
rect 104 43420 1916 43488
rect 104 43364 114 43420
rect 170 43364 238 43420
rect 294 43364 362 43420
rect 418 43364 486 43420
rect 542 43364 610 43420
rect 666 43364 734 43420
rect 790 43364 858 43420
rect 914 43364 982 43420
rect 1038 43364 1106 43420
rect 1162 43364 1230 43420
rect 1286 43364 1354 43420
rect 1410 43364 1478 43420
rect 1534 43364 1602 43420
rect 1658 43364 1726 43420
rect 1782 43364 1850 43420
rect 1906 43364 1916 43420
rect 104 43296 1916 43364
rect 104 43240 114 43296
rect 170 43240 238 43296
rect 294 43240 362 43296
rect 418 43240 486 43296
rect 542 43240 610 43296
rect 666 43240 734 43296
rect 790 43240 858 43296
rect 914 43240 982 43296
rect 1038 43240 1106 43296
rect 1162 43240 1230 43296
rect 1286 43240 1354 43296
rect 1410 43240 1478 43296
rect 1534 43240 1602 43296
rect 1658 43240 1726 43296
rect 1782 43240 1850 43296
rect 1906 43240 1916 43296
rect 104 43172 1916 43240
rect 104 43116 114 43172
rect 170 43116 238 43172
rect 294 43116 362 43172
rect 418 43116 486 43172
rect 542 43116 610 43172
rect 666 43116 734 43172
rect 790 43116 858 43172
rect 914 43116 982 43172
rect 1038 43116 1106 43172
rect 1162 43116 1230 43172
rect 1286 43116 1354 43172
rect 1410 43116 1478 43172
rect 1534 43116 1602 43172
rect 1658 43116 1726 43172
rect 1782 43116 1850 43172
rect 1906 43116 1916 43172
rect 104 43048 1916 43116
rect 104 42992 114 43048
rect 170 42992 238 43048
rect 294 42992 362 43048
rect 418 42992 486 43048
rect 542 42992 610 43048
rect 666 42992 734 43048
rect 790 42992 858 43048
rect 914 42992 982 43048
rect 1038 42992 1106 43048
rect 1162 42992 1230 43048
rect 1286 42992 1354 43048
rect 1410 42992 1478 43048
rect 1534 42992 1602 43048
rect 1658 42992 1726 43048
rect 1782 42992 1850 43048
rect 1906 42992 1916 43048
rect 104 42982 1916 42992
rect 104 42487 1916 42497
rect 104 42431 114 42487
rect 170 42431 238 42487
rect 294 42431 362 42487
rect 418 42431 486 42487
rect 542 42431 610 42487
rect 666 42431 734 42487
rect 790 42431 858 42487
rect 914 42431 982 42487
rect 1038 42431 1106 42487
rect 1162 42431 1230 42487
rect 1286 42431 1354 42487
rect 1410 42431 1478 42487
rect 1534 42431 1602 42487
rect 1658 42431 1726 42487
rect 1782 42431 1850 42487
rect 1906 42431 1916 42487
rect 104 42363 1916 42431
rect 104 42307 114 42363
rect 170 42307 238 42363
rect 294 42307 362 42363
rect 418 42307 486 42363
rect 542 42307 610 42363
rect 666 42307 734 42363
rect 790 42307 858 42363
rect 914 42307 982 42363
rect 1038 42307 1106 42363
rect 1162 42307 1230 42363
rect 1286 42307 1354 42363
rect 1410 42307 1478 42363
rect 1534 42307 1602 42363
rect 1658 42307 1726 42363
rect 1782 42307 1850 42363
rect 1906 42307 1916 42363
rect 104 42239 1916 42307
rect 104 42183 114 42239
rect 170 42183 238 42239
rect 294 42183 362 42239
rect 418 42183 486 42239
rect 542 42183 610 42239
rect 666 42183 734 42239
rect 790 42183 858 42239
rect 914 42183 982 42239
rect 1038 42183 1106 42239
rect 1162 42183 1230 42239
rect 1286 42183 1354 42239
rect 1410 42183 1478 42239
rect 1534 42183 1602 42239
rect 1658 42183 1726 42239
rect 1782 42183 1850 42239
rect 1906 42183 1916 42239
rect 104 42115 1916 42183
rect 104 42059 114 42115
rect 170 42059 238 42115
rect 294 42059 362 42115
rect 418 42059 486 42115
rect 542 42059 610 42115
rect 666 42059 734 42115
rect 790 42059 858 42115
rect 914 42059 982 42115
rect 1038 42059 1106 42115
rect 1162 42059 1230 42115
rect 1286 42059 1354 42115
rect 1410 42059 1478 42115
rect 1534 42059 1602 42115
rect 1658 42059 1726 42115
rect 1782 42059 1850 42115
rect 1906 42059 1916 42115
rect 104 41991 1916 42059
rect 104 41935 114 41991
rect 170 41935 238 41991
rect 294 41935 362 41991
rect 418 41935 486 41991
rect 542 41935 610 41991
rect 666 41935 734 41991
rect 790 41935 858 41991
rect 914 41935 982 41991
rect 1038 41935 1106 41991
rect 1162 41935 1230 41991
rect 1286 41935 1354 41991
rect 1410 41935 1478 41991
rect 1534 41935 1602 41991
rect 1658 41935 1726 41991
rect 1782 41935 1850 41991
rect 1906 41935 1916 41991
rect 104 41867 1916 41935
rect 104 41811 114 41867
rect 170 41811 238 41867
rect 294 41811 362 41867
rect 418 41811 486 41867
rect 542 41811 610 41867
rect 666 41811 734 41867
rect 790 41811 858 41867
rect 914 41811 982 41867
rect 1038 41811 1106 41867
rect 1162 41811 1230 41867
rect 1286 41811 1354 41867
rect 1410 41811 1478 41867
rect 1534 41811 1602 41867
rect 1658 41811 1726 41867
rect 1782 41811 1850 41867
rect 1906 41811 1916 41867
rect 104 41743 1916 41811
rect 104 41687 114 41743
rect 170 41687 238 41743
rect 294 41687 362 41743
rect 418 41687 486 41743
rect 542 41687 610 41743
rect 666 41687 734 41743
rect 790 41687 858 41743
rect 914 41687 982 41743
rect 1038 41687 1106 41743
rect 1162 41687 1230 41743
rect 1286 41687 1354 41743
rect 1410 41687 1478 41743
rect 1534 41687 1602 41743
rect 1658 41687 1726 41743
rect 1782 41687 1850 41743
rect 1906 41687 1916 41743
rect 104 41619 1916 41687
rect 104 41563 114 41619
rect 170 41563 238 41619
rect 294 41563 362 41619
rect 418 41563 486 41619
rect 542 41563 610 41619
rect 666 41563 734 41619
rect 790 41563 858 41619
rect 914 41563 982 41619
rect 1038 41563 1106 41619
rect 1162 41563 1230 41619
rect 1286 41563 1354 41619
rect 1410 41563 1478 41619
rect 1534 41563 1602 41619
rect 1658 41563 1726 41619
rect 1782 41563 1850 41619
rect 1906 41563 1916 41619
rect 104 41495 1916 41563
rect 104 41439 114 41495
rect 170 41439 238 41495
rect 294 41439 362 41495
rect 418 41439 486 41495
rect 542 41439 610 41495
rect 666 41439 734 41495
rect 790 41439 858 41495
rect 914 41439 982 41495
rect 1038 41439 1106 41495
rect 1162 41439 1230 41495
rect 1286 41439 1354 41495
rect 1410 41439 1478 41495
rect 1534 41439 1602 41495
rect 1658 41439 1726 41495
rect 1782 41439 1850 41495
rect 1906 41439 1916 41495
rect 104 41371 1916 41439
rect 104 41315 114 41371
rect 170 41315 238 41371
rect 294 41315 362 41371
rect 418 41315 486 41371
rect 542 41315 610 41371
rect 666 41315 734 41371
rect 790 41315 858 41371
rect 914 41315 982 41371
rect 1038 41315 1106 41371
rect 1162 41315 1230 41371
rect 1286 41315 1354 41371
rect 1410 41315 1478 41371
rect 1534 41315 1602 41371
rect 1658 41315 1726 41371
rect 1782 41315 1850 41371
rect 1906 41315 1916 41371
rect 104 41305 1916 41315
rect 104 40891 1916 40901
rect 104 40835 114 40891
rect 170 40835 238 40891
rect 294 40835 362 40891
rect 418 40835 486 40891
rect 542 40835 610 40891
rect 666 40835 734 40891
rect 790 40835 858 40891
rect 914 40835 982 40891
rect 1038 40835 1106 40891
rect 1162 40835 1230 40891
rect 1286 40835 1354 40891
rect 1410 40835 1478 40891
rect 1534 40835 1602 40891
rect 1658 40835 1726 40891
rect 1782 40835 1850 40891
rect 1906 40835 1916 40891
rect 104 40767 1916 40835
rect 104 40711 114 40767
rect 170 40711 238 40767
rect 294 40711 362 40767
rect 418 40711 486 40767
rect 542 40711 610 40767
rect 666 40711 734 40767
rect 790 40711 858 40767
rect 914 40711 982 40767
rect 1038 40711 1106 40767
rect 1162 40711 1230 40767
rect 1286 40711 1354 40767
rect 1410 40711 1478 40767
rect 1534 40711 1602 40767
rect 1658 40711 1726 40767
rect 1782 40711 1850 40767
rect 1906 40711 1916 40767
rect 104 40643 1916 40711
rect 104 40587 114 40643
rect 170 40587 238 40643
rect 294 40587 362 40643
rect 418 40587 486 40643
rect 542 40587 610 40643
rect 666 40587 734 40643
rect 790 40587 858 40643
rect 914 40587 982 40643
rect 1038 40587 1106 40643
rect 1162 40587 1230 40643
rect 1286 40587 1354 40643
rect 1410 40587 1478 40643
rect 1534 40587 1602 40643
rect 1658 40587 1726 40643
rect 1782 40587 1850 40643
rect 1906 40587 1916 40643
rect 104 40519 1916 40587
rect 104 40463 114 40519
rect 170 40463 238 40519
rect 294 40463 362 40519
rect 418 40463 486 40519
rect 542 40463 610 40519
rect 666 40463 734 40519
rect 790 40463 858 40519
rect 914 40463 982 40519
rect 1038 40463 1106 40519
rect 1162 40463 1230 40519
rect 1286 40463 1354 40519
rect 1410 40463 1478 40519
rect 1534 40463 1602 40519
rect 1658 40463 1726 40519
rect 1782 40463 1850 40519
rect 1906 40463 1916 40519
rect 104 40395 1916 40463
rect 104 40339 114 40395
rect 170 40339 238 40395
rect 294 40339 362 40395
rect 418 40339 486 40395
rect 542 40339 610 40395
rect 666 40339 734 40395
rect 790 40339 858 40395
rect 914 40339 982 40395
rect 1038 40339 1106 40395
rect 1162 40339 1230 40395
rect 1286 40339 1354 40395
rect 1410 40339 1478 40395
rect 1534 40339 1602 40395
rect 1658 40339 1726 40395
rect 1782 40339 1850 40395
rect 1906 40339 1916 40395
rect 104 40271 1916 40339
rect 104 40215 114 40271
rect 170 40215 238 40271
rect 294 40215 362 40271
rect 418 40215 486 40271
rect 542 40215 610 40271
rect 666 40215 734 40271
rect 790 40215 858 40271
rect 914 40215 982 40271
rect 1038 40215 1106 40271
rect 1162 40215 1230 40271
rect 1286 40215 1354 40271
rect 1410 40215 1478 40271
rect 1534 40215 1602 40271
rect 1658 40215 1726 40271
rect 1782 40215 1850 40271
rect 1906 40215 1916 40271
rect 104 40147 1916 40215
rect 104 40091 114 40147
rect 170 40091 238 40147
rect 294 40091 362 40147
rect 418 40091 486 40147
rect 542 40091 610 40147
rect 666 40091 734 40147
rect 790 40091 858 40147
rect 914 40091 982 40147
rect 1038 40091 1106 40147
rect 1162 40091 1230 40147
rect 1286 40091 1354 40147
rect 1410 40091 1478 40147
rect 1534 40091 1602 40147
rect 1658 40091 1726 40147
rect 1782 40091 1850 40147
rect 1906 40091 1916 40147
rect 104 40023 1916 40091
rect 104 39967 114 40023
rect 170 39967 238 40023
rect 294 39967 362 40023
rect 418 39967 486 40023
rect 542 39967 610 40023
rect 666 39967 734 40023
rect 790 39967 858 40023
rect 914 39967 982 40023
rect 1038 39967 1106 40023
rect 1162 39967 1230 40023
rect 1286 39967 1354 40023
rect 1410 39967 1478 40023
rect 1534 39967 1602 40023
rect 1658 39967 1726 40023
rect 1782 39967 1850 40023
rect 1906 39967 1916 40023
rect 104 39899 1916 39967
rect 104 39843 114 39899
rect 170 39843 238 39899
rect 294 39843 362 39899
rect 418 39843 486 39899
rect 542 39843 610 39899
rect 666 39843 734 39899
rect 790 39843 858 39899
rect 914 39843 982 39899
rect 1038 39843 1106 39899
rect 1162 39843 1230 39899
rect 1286 39843 1354 39899
rect 1410 39843 1478 39899
rect 1534 39843 1602 39899
rect 1658 39843 1726 39899
rect 1782 39843 1850 39899
rect 1906 39843 1916 39899
rect 104 39775 1916 39843
rect 104 39719 114 39775
rect 170 39719 238 39775
rect 294 39719 362 39775
rect 418 39719 486 39775
rect 542 39719 610 39775
rect 666 39719 734 39775
rect 790 39719 858 39775
rect 914 39719 982 39775
rect 1038 39719 1106 39775
rect 1162 39719 1230 39775
rect 1286 39719 1354 39775
rect 1410 39719 1478 39775
rect 1534 39719 1602 39775
rect 1658 39719 1726 39775
rect 1782 39719 1850 39775
rect 1906 39719 1916 39775
rect 104 39709 1916 39719
rect 104 39244 1916 39254
rect 104 39188 114 39244
rect 170 39188 238 39244
rect 294 39188 362 39244
rect 418 39188 486 39244
rect 542 39188 610 39244
rect 666 39188 734 39244
rect 790 39188 858 39244
rect 914 39188 982 39244
rect 1038 39188 1106 39244
rect 1162 39188 1230 39244
rect 1286 39188 1354 39244
rect 1410 39188 1478 39244
rect 1534 39188 1602 39244
rect 1658 39188 1726 39244
rect 1782 39188 1850 39244
rect 1906 39188 1916 39244
rect 104 39120 1916 39188
rect 104 39064 114 39120
rect 170 39064 238 39120
rect 294 39064 362 39120
rect 418 39064 486 39120
rect 542 39064 610 39120
rect 666 39064 734 39120
rect 790 39064 858 39120
rect 914 39064 982 39120
rect 1038 39064 1106 39120
rect 1162 39064 1230 39120
rect 1286 39064 1354 39120
rect 1410 39064 1478 39120
rect 1534 39064 1602 39120
rect 1658 39064 1726 39120
rect 1782 39064 1850 39120
rect 1906 39064 1916 39120
rect 104 38996 1916 39064
rect 104 38940 114 38996
rect 170 38940 238 38996
rect 294 38940 362 38996
rect 418 38940 486 38996
rect 542 38940 610 38996
rect 666 38940 734 38996
rect 790 38940 858 38996
rect 914 38940 982 38996
rect 1038 38940 1106 38996
rect 1162 38940 1230 38996
rect 1286 38940 1354 38996
rect 1410 38940 1478 38996
rect 1534 38940 1602 38996
rect 1658 38940 1726 38996
rect 1782 38940 1850 38996
rect 1906 38940 1916 38996
rect 104 38872 1916 38940
rect 104 38816 114 38872
rect 170 38816 238 38872
rect 294 38816 362 38872
rect 418 38816 486 38872
rect 542 38816 610 38872
rect 666 38816 734 38872
rect 790 38816 858 38872
rect 914 38816 982 38872
rect 1038 38816 1106 38872
rect 1162 38816 1230 38872
rect 1286 38816 1354 38872
rect 1410 38816 1478 38872
rect 1534 38816 1602 38872
rect 1658 38816 1726 38872
rect 1782 38816 1850 38872
rect 1906 38816 1916 38872
rect 104 38748 1916 38816
rect 104 38692 114 38748
rect 170 38692 238 38748
rect 294 38692 362 38748
rect 418 38692 486 38748
rect 542 38692 610 38748
rect 666 38692 734 38748
rect 790 38692 858 38748
rect 914 38692 982 38748
rect 1038 38692 1106 38748
rect 1162 38692 1230 38748
rect 1286 38692 1354 38748
rect 1410 38692 1478 38748
rect 1534 38692 1602 38748
rect 1658 38692 1726 38748
rect 1782 38692 1850 38748
rect 1906 38692 1916 38748
rect 104 38624 1916 38692
rect 104 38568 114 38624
rect 170 38568 238 38624
rect 294 38568 362 38624
rect 418 38568 486 38624
rect 542 38568 610 38624
rect 666 38568 734 38624
rect 790 38568 858 38624
rect 914 38568 982 38624
rect 1038 38568 1106 38624
rect 1162 38568 1230 38624
rect 1286 38568 1354 38624
rect 1410 38568 1478 38624
rect 1534 38568 1602 38624
rect 1658 38568 1726 38624
rect 1782 38568 1850 38624
rect 1906 38568 1916 38624
rect 104 38500 1916 38568
rect 104 38444 114 38500
rect 170 38444 238 38500
rect 294 38444 362 38500
rect 418 38444 486 38500
rect 542 38444 610 38500
rect 666 38444 734 38500
rect 790 38444 858 38500
rect 914 38444 982 38500
rect 1038 38444 1106 38500
rect 1162 38444 1230 38500
rect 1286 38444 1354 38500
rect 1410 38444 1478 38500
rect 1534 38444 1602 38500
rect 1658 38444 1726 38500
rect 1782 38444 1850 38500
rect 1906 38444 1916 38500
rect 104 38376 1916 38444
rect 104 38320 114 38376
rect 170 38320 238 38376
rect 294 38320 362 38376
rect 418 38320 486 38376
rect 542 38320 610 38376
rect 666 38320 734 38376
rect 790 38320 858 38376
rect 914 38320 982 38376
rect 1038 38320 1106 38376
rect 1162 38320 1230 38376
rect 1286 38320 1354 38376
rect 1410 38320 1478 38376
rect 1534 38320 1602 38376
rect 1658 38320 1726 38376
rect 1782 38320 1850 38376
rect 1906 38320 1916 38376
rect 104 38252 1916 38320
rect 104 38196 114 38252
rect 170 38196 238 38252
rect 294 38196 362 38252
rect 418 38196 486 38252
rect 542 38196 610 38252
rect 666 38196 734 38252
rect 790 38196 858 38252
rect 914 38196 982 38252
rect 1038 38196 1106 38252
rect 1162 38196 1230 38252
rect 1286 38196 1354 38252
rect 1410 38196 1478 38252
rect 1534 38196 1602 38252
rect 1658 38196 1726 38252
rect 1782 38196 1850 38252
rect 1906 38196 1916 38252
rect 104 38128 1916 38196
rect 104 38072 114 38128
rect 170 38072 238 38128
rect 294 38072 362 38128
rect 418 38072 486 38128
rect 542 38072 610 38128
rect 666 38072 734 38128
rect 790 38072 858 38128
rect 914 38072 982 38128
rect 1038 38072 1106 38128
rect 1162 38072 1230 38128
rect 1286 38072 1354 38128
rect 1410 38072 1478 38128
rect 1534 38072 1602 38128
rect 1658 38072 1726 38128
rect 1782 38072 1850 38128
rect 1906 38072 1916 38128
rect 104 38004 1916 38072
rect 104 37948 114 38004
rect 170 37948 238 38004
rect 294 37948 362 38004
rect 418 37948 486 38004
rect 542 37948 610 38004
rect 666 37948 734 38004
rect 790 37948 858 38004
rect 914 37948 982 38004
rect 1038 37948 1106 38004
rect 1162 37948 1230 38004
rect 1286 37948 1354 38004
rect 1410 37948 1478 38004
rect 1534 37948 1602 38004
rect 1658 37948 1726 38004
rect 1782 37948 1850 38004
rect 1906 37948 1916 38004
rect 104 37880 1916 37948
rect 104 37824 114 37880
rect 170 37824 238 37880
rect 294 37824 362 37880
rect 418 37824 486 37880
rect 542 37824 610 37880
rect 666 37824 734 37880
rect 790 37824 858 37880
rect 914 37824 982 37880
rect 1038 37824 1106 37880
rect 1162 37824 1230 37880
rect 1286 37824 1354 37880
rect 1410 37824 1478 37880
rect 1534 37824 1602 37880
rect 1658 37824 1726 37880
rect 1782 37824 1850 37880
rect 1906 37824 1916 37880
rect 104 37756 1916 37824
rect 104 37700 114 37756
rect 170 37700 238 37756
rect 294 37700 362 37756
rect 418 37700 486 37756
rect 542 37700 610 37756
rect 666 37700 734 37756
rect 790 37700 858 37756
rect 914 37700 982 37756
rect 1038 37700 1106 37756
rect 1162 37700 1230 37756
rect 1286 37700 1354 37756
rect 1410 37700 1478 37756
rect 1534 37700 1602 37756
rect 1658 37700 1726 37756
rect 1782 37700 1850 37756
rect 1906 37700 1916 37756
rect 104 37632 1916 37700
rect 104 37576 114 37632
rect 170 37576 238 37632
rect 294 37576 362 37632
rect 418 37576 486 37632
rect 542 37576 610 37632
rect 666 37576 734 37632
rect 790 37576 858 37632
rect 914 37576 982 37632
rect 1038 37576 1106 37632
rect 1162 37576 1230 37632
rect 1286 37576 1354 37632
rect 1410 37576 1478 37632
rect 1534 37576 1602 37632
rect 1658 37576 1726 37632
rect 1782 37576 1850 37632
rect 1906 37576 1916 37632
rect 104 37508 1916 37576
rect 104 37452 114 37508
rect 170 37452 238 37508
rect 294 37452 362 37508
rect 418 37452 486 37508
rect 542 37452 610 37508
rect 666 37452 734 37508
rect 790 37452 858 37508
rect 914 37452 982 37508
rect 1038 37452 1106 37508
rect 1162 37452 1230 37508
rect 1286 37452 1354 37508
rect 1410 37452 1478 37508
rect 1534 37452 1602 37508
rect 1658 37452 1726 37508
rect 1782 37452 1850 37508
rect 1906 37452 1916 37508
rect 104 37384 1916 37452
rect 104 37328 114 37384
rect 170 37328 238 37384
rect 294 37328 362 37384
rect 418 37328 486 37384
rect 542 37328 610 37384
rect 666 37328 734 37384
rect 790 37328 858 37384
rect 914 37328 982 37384
rect 1038 37328 1106 37384
rect 1162 37328 1230 37384
rect 1286 37328 1354 37384
rect 1410 37328 1478 37384
rect 1534 37328 1602 37384
rect 1658 37328 1726 37384
rect 1782 37328 1850 37384
rect 1906 37328 1916 37384
rect 104 37260 1916 37328
rect 104 37204 114 37260
rect 170 37204 238 37260
rect 294 37204 362 37260
rect 418 37204 486 37260
rect 542 37204 610 37260
rect 666 37204 734 37260
rect 790 37204 858 37260
rect 914 37204 982 37260
rect 1038 37204 1106 37260
rect 1162 37204 1230 37260
rect 1286 37204 1354 37260
rect 1410 37204 1478 37260
rect 1534 37204 1602 37260
rect 1658 37204 1726 37260
rect 1782 37204 1850 37260
rect 1906 37204 1916 37260
rect 104 37136 1916 37204
rect 104 37080 114 37136
rect 170 37080 238 37136
rect 294 37080 362 37136
rect 418 37080 486 37136
rect 542 37080 610 37136
rect 666 37080 734 37136
rect 790 37080 858 37136
rect 914 37080 982 37136
rect 1038 37080 1106 37136
rect 1162 37080 1230 37136
rect 1286 37080 1354 37136
rect 1410 37080 1478 37136
rect 1534 37080 1602 37136
rect 1658 37080 1726 37136
rect 1782 37080 1850 37136
rect 1906 37080 1916 37136
rect 104 37012 1916 37080
rect 104 36956 114 37012
rect 170 36956 238 37012
rect 294 36956 362 37012
rect 418 36956 486 37012
rect 542 36956 610 37012
rect 666 36956 734 37012
rect 790 36956 858 37012
rect 914 36956 982 37012
rect 1038 36956 1106 37012
rect 1162 36956 1230 37012
rect 1286 36956 1354 37012
rect 1410 36956 1478 37012
rect 1534 36956 1602 37012
rect 1658 36956 1726 37012
rect 1782 36956 1850 37012
rect 1906 36956 1916 37012
rect 104 36888 1916 36956
rect 104 36832 114 36888
rect 170 36832 238 36888
rect 294 36832 362 36888
rect 418 36832 486 36888
rect 542 36832 610 36888
rect 666 36832 734 36888
rect 790 36832 858 36888
rect 914 36832 982 36888
rect 1038 36832 1106 36888
rect 1162 36832 1230 36888
rect 1286 36832 1354 36888
rect 1410 36832 1478 36888
rect 1534 36832 1602 36888
rect 1658 36832 1726 36888
rect 1782 36832 1850 36888
rect 1906 36832 1916 36888
rect 104 36764 1916 36832
rect 104 36708 114 36764
rect 170 36708 238 36764
rect 294 36708 362 36764
rect 418 36708 486 36764
rect 542 36708 610 36764
rect 666 36708 734 36764
rect 790 36708 858 36764
rect 914 36708 982 36764
rect 1038 36708 1106 36764
rect 1162 36708 1230 36764
rect 1286 36708 1354 36764
rect 1410 36708 1478 36764
rect 1534 36708 1602 36764
rect 1658 36708 1726 36764
rect 1782 36708 1850 36764
rect 1906 36708 1916 36764
rect 104 36640 1916 36708
rect 104 36584 114 36640
rect 170 36584 238 36640
rect 294 36584 362 36640
rect 418 36584 486 36640
rect 542 36584 610 36640
rect 666 36584 734 36640
rect 790 36584 858 36640
rect 914 36584 982 36640
rect 1038 36584 1106 36640
rect 1162 36584 1230 36640
rect 1286 36584 1354 36640
rect 1410 36584 1478 36640
rect 1534 36584 1602 36640
rect 1658 36584 1726 36640
rect 1782 36584 1850 36640
rect 1906 36584 1916 36640
rect 104 36574 1916 36584
rect 104 36059 1916 36069
rect 104 36003 114 36059
rect 170 36003 238 36059
rect 294 36003 362 36059
rect 418 36003 486 36059
rect 542 36003 610 36059
rect 666 36003 734 36059
rect 790 36003 858 36059
rect 914 36003 982 36059
rect 1038 36003 1106 36059
rect 1162 36003 1230 36059
rect 1286 36003 1354 36059
rect 1410 36003 1478 36059
rect 1534 36003 1602 36059
rect 1658 36003 1726 36059
rect 1782 36003 1850 36059
rect 1906 36003 1916 36059
rect 104 35935 1916 36003
rect 104 35879 114 35935
rect 170 35879 238 35935
rect 294 35879 362 35935
rect 418 35879 486 35935
rect 542 35879 610 35935
rect 666 35879 734 35935
rect 790 35879 858 35935
rect 914 35879 982 35935
rect 1038 35879 1106 35935
rect 1162 35879 1230 35935
rect 1286 35879 1354 35935
rect 1410 35879 1478 35935
rect 1534 35879 1602 35935
rect 1658 35879 1726 35935
rect 1782 35879 1850 35935
rect 1906 35879 1916 35935
rect 104 35811 1916 35879
rect 104 35755 114 35811
rect 170 35755 238 35811
rect 294 35755 362 35811
rect 418 35755 486 35811
rect 542 35755 610 35811
rect 666 35755 734 35811
rect 790 35755 858 35811
rect 914 35755 982 35811
rect 1038 35755 1106 35811
rect 1162 35755 1230 35811
rect 1286 35755 1354 35811
rect 1410 35755 1478 35811
rect 1534 35755 1602 35811
rect 1658 35755 1726 35811
rect 1782 35755 1850 35811
rect 1906 35755 1916 35811
rect 104 35687 1916 35755
rect 104 35631 114 35687
rect 170 35631 238 35687
rect 294 35631 362 35687
rect 418 35631 486 35687
rect 542 35631 610 35687
rect 666 35631 734 35687
rect 790 35631 858 35687
rect 914 35631 982 35687
rect 1038 35631 1106 35687
rect 1162 35631 1230 35687
rect 1286 35631 1354 35687
rect 1410 35631 1478 35687
rect 1534 35631 1602 35687
rect 1658 35631 1726 35687
rect 1782 35631 1850 35687
rect 1906 35631 1916 35687
rect 104 35563 1916 35631
rect 104 35507 114 35563
rect 170 35507 238 35563
rect 294 35507 362 35563
rect 418 35507 486 35563
rect 542 35507 610 35563
rect 666 35507 734 35563
rect 790 35507 858 35563
rect 914 35507 982 35563
rect 1038 35507 1106 35563
rect 1162 35507 1230 35563
rect 1286 35507 1354 35563
rect 1410 35507 1478 35563
rect 1534 35507 1602 35563
rect 1658 35507 1726 35563
rect 1782 35507 1850 35563
rect 1906 35507 1916 35563
rect 104 35439 1916 35507
rect 104 35383 114 35439
rect 170 35383 238 35439
rect 294 35383 362 35439
rect 418 35383 486 35439
rect 542 35383 610 35439
rect 666 35383 734 35439
rect 790 35383 858 35439
rect 914 35383 982 35439
rect 1038 35383 1106 35439
rect 1162 35383 1230 35439
rect 1286 35383 1354 35439
rect 1410 35383 1478 35439
rect 1534 35383 1602 35439
rect 1658 35383 1726 35439
rect 1782 35383 1850 35439
rect 1906 35383 1916 35439
rect 104 35315 1916 35383
rect 104 35259 114 35315
rect 170 35259 238 35315
rect 294 35259 362 35315
rect 418 35259 486 35315
rect 542 35259 610 35315
rect 666 35259 734 35315
rect 790 35259 858 35315
rect 914 35259 982 35315
rect 1038 35259 1106 35315
rect 1162 35259 1230 35315
rect 1286 35259 1354 35315
rect 1410 35259 1478 35315
rect 1534 35259 1602 35315
rect 1658 35259 1726 35315
rect 1782 35259 1850 35315
rect 1906 35259 1916 35315
rect 104 35191 1916 35259
rect 104 35135 114 35191
rect 170 35135 238 35191
rect 294 35135 362 35191
rect 418 35135 486 35191
rect 542 35135 610 35191
rect 666 35135 734 35191
rect 790 35135 858 35191
rect 914 35135 982 35191
rect 1038 35135 1106 35191
rect 1162 35135 1230 35191
rect 1286 35135 1354 35191
rect 1410 35135 1478 35191
rect 1534 35135 1602 35191
rect 1658 35135 1726 35191
rect 1782 35135 1850 35191
rect 1906 35135 1916 35191
rect 104 35067 1916 35135
rect 104 35011 114 35067
rect 170 35011 238 35067
rect 294 35011 362 35067
rect 418 35011 486 35067
rect 542 35011 610 35067
rect 666 35011 734 35067
rect 790 35011 858 35067
rect 914 35011 982 35067
rect 1038 35011 1106 35067
rect 1162 35011 1230 35067
rect 1286 35011 1354 35067
rect 1410 35011 1478 35067
rect 1534 35011 1602 35067
rect 1658 35011 1726 35067
rect 1782 35011 1850 35067
rect 1906 35011 1916 35067
rect 104 34943 1916 35011
rect 104 34887 114 34943
rect 170 34887 238 34943
rect 294 34887 362 34943
rect 418 34887 486 34943
rect 542 34887 610 34943
rect 666 34887 734 34943
rect 790 34887 858 34943
rect 914 34887 982 34943
rect 1038 34887 1106 34943
rect 1162 34887 1230 34943
rect 1286 34887 1354 34943
rect 1410 34887 1478 34943
rect 1534 34887 1602 34943
rect 1658 34887 1726 34943
rect 1782 34887 1850 34943
rect 1906 34887 1916 34943
rect 104 34819 1916 34887
rect 104 34763 114 34819
rect 170 34763 238 34819
rect 294 34763 362 34819
rect 418 34763 486 34819
rect 542 34763 610 34819
rect 666 34763 734 34819
rect 790 34763 858 34819
rect 914 34763 982 34819
rect 1038 34763 1106 34819
rect 1162 34763 1230 34819
rect 1286 34763 1354 34819
rect 1410 34763 1478 34819
rect 1534 34763 1602 34819
rect 1658 34763 1726 34819
rect 1782 34763 1850 34819
rect 1906 34763 1916 34819
rect 104 34695 1916 34763
rect 104 34639 114 34695
rect 170 34639 238 34695
rect 294 34639 362 34695
rect 418 34639 486 34695
rect 542 34639 610 34695
rect 666 34639 734 34695
rect 790 34639 858 34695
rect 914 34639 982 34695
rect 1038 34639 1106 34695
rect 1162 34639 1230 34695
rect 1286 34639 1354 34695
rect 1410 34639 1478 34695
rect 1534 34639 1602 34695
rect 1658 34639 1726 34695
rect 1782 34639 1850 34695
rect 1906 34639 1916 34695
rect 104 34571 1916 34639
rect 104 34515 114 34571
rect 170 34515 238 34571
rect 294 34515 362 34571
rect 418 34515 486 34571
rect 542 34515 610 34571
rect 666 34515 734 34571
rect 790 34515 858 34571
rect 914 34515 982 34571
rect 1038 34515 1106 34571
rect 1162 34515 1230 34571
rect 1286 34515 1354 34571
rect 1410 34515 1478 34571
rect 1534 34515 1602 34571
rect 1658 34515 1726 34571
rect 1782 34515 1850 34571
rect 1906 34515 1916 34571
rect 104 34447 1916 34515
rect 104 34391 114 34447
rect 170 34391 238 34447
rect 294 34391 362 34447
rect 418 34391 486 34447
rect 542 34391 610 34447
rect 666 34391 734 34447
rect 790 34391 858 34447
rect 914 34391 982 34447
rect 1038 34391 1106 34447
rect 1162 34391 1230 34447
rect 1286 34391 1354 34447
rect 1410 34391 1478 34447
rect 1534 34391 1602 34447
rect 1658 34391 1726 34447
rect 1782 34391 1850 34447
rect 1906 34391 1916 34447
rect 104 34323 1916 34391
rect 104 34267 114 34323
rect 170 34267 238 34323
rect 294 34267 362 34323
rect 418 34267 486 34323
rect 542 34267 610 34323
rect 666 34267 734 34323
rect 790 34267 858 34323
rect 914 34267 982 34323
rect 1038 34267 1106 34323
rect 1162 34267 1230 34323
rect 1286 34267 1354 34323
rect 1410 34267 1478 34323
rect 1534 34267 1602 34323
rect 1658 34267 1726 34323
rect 1782 34267 1850 34323
rect 1906 34267 1916 34323
rect 104 34199 1916 34267
rect 104 34143 114 34199
rect 170 34143 238 34199
rect 294 34143 362 34199
rect 418 34143 486 34199
rect 542 34143 610 34199
rect 666 34143 734 34199
rect 790 34143 858 34199
rect 914 34143 982 34199
rect 1038 34143 1106 34199
rect 1162 34143 1230 34199
rect 1286 34143 1354 34199
rect 1410 34143 1478 34199
rect 1534 34143 1602 34199
rect 1658 34143 1726 34199
rect 1782 34143 1850 34199
rect 1906 34143 1916 34199
rect 104 34075 1916 34143
rect 104 34019 114 34075
rect 170 34019 238 34075
rect 294 34019 362 34075
rect 418 34019 486 34075
rect 542 34019 610 34075
rect 666 34019 734 34075
rect 790 34019 858 34075
rect 914 34019 982 34075
rect 1038 34019 1106 34075
rect 1162 34019 1230 34075
rect 1286 34019 1354 34075
rect 1410 34019 1478 34075
rect 1534 34019 1602 34075
rect 1658 34019 1726 34075
rect 1782 34019 1850 34075
rect 1906 34019 1916 34075
rect 104 33951 1916 34019
rect 104 33895 114 33951
rect 170 33895 238 33951
rect 294 33895 362 33951
rect 418 33895 486 33951
rect 542 33895 610 33951
rect 666 33895 734 33951
rect 790 33895 858 33951
rect 914 33895 982 33951
rect 1038 33895 1106 33951
rect 1162 33895 1230 33951
rect 1286 33895 1354 33951
rect 1410 33895 1478 33951
rect 1534 33895 1602 33951
rect 1658 33895 1726 33951
rect 1782 33895 1850 33951
rect 1906 33895 1916 33951
rect 104 33827 1916 33895
rect 104 33771 114 33827
rect 170 33771 238 33827
rect 294 33771 362 33827
rect 418 33771 486 33827
rect 542 33771 610 33827
rect 666 33771 734 33827
rect 790 33771 858 33827
rect 914 33771 982 33827
rect 1038 33771 1106 33827
rect 1162 33771 1230 33827
rect 1286 33771 1354 33827
rect 1410 33771 1478 33827
rect 1534 33771 1602 33827
rect 1658 33771 1726 33827
rect 1782 33771 1850 33827
rect 1906 33771 1916 33827
rect 104 33703 1916 33771
rect 104 33647 114 33703
rect 170 33647 238 33703
rect 294 33647 362 33703
rect 418 33647 486 33703
rect 542 33647 610 33703
rect 666 33647 734 33703
rect 790 33647 858 33703
rect 914 33647 982 33703
rect 1038 33647 1106 33703
rect 1162 33647 1230 33703
rect 1286 33647 1354 33703
rect 1410 33647 1478 33703
rect 1534 33647 1602 33703
rect 1658 33647 1726 33703
rect 1782 33647 1850 33703
rect 1906 33647 1916 33703
rect 104 33579 1916 33647
rect 104 33523 114 33579
rect 170 33523 238 33579
rect 294 33523 362 33579
rect 418 33523 486 33579
rect 542 33523 610 33579
rect 666 33523 734 33579
rect 790 33523 858 33579
rect 914 33523 982 33579
rect 1038 33523 1106 33579
rect 1162 33523 1230 33579
rect 1286 33523 1354 33579
rect 1410 33523 1478 33579
rect 1534 33523 1602 33579
rect 1658 33523 1726 33579
rect 1782 33523 1850 33579
rect 1906 33523 1916 33579
rect 104 33455 1916 33523
rect 104 33399 114 33455
rect 170 33399 238 33455
rect 294 33399 362 33455
rect 418 33399 486 33455
rect 542 33399 610 33455
rect 666 33399 734 33455
rect 790 33399 858 33455
rect 914 33399 982 33455
rect 1038 33399 1106 33455
rect 1162 33399 1230 33455
rect 1286 33399 1354 33455
rect 1410 33399 1478 33455
rect 1534 33399 1602 33455
rect 1658 33399 1726 33455
rect 1782 33399 1850 33455
rect 1906 33399 1916 33455
rect 104 33389 1916 33399
rect 104 32844 1916 32854
rect 104 32788 114 32844
rect 170 32788 238 32844
rect 294 32788 362 32844
rect 418 32788 486 32844
rect 542 32788 610 32844
rect 666 32788 734 32844
rect 790 32788 858 32844
rect 914 32788 982 32844
rect 1038 32788 1106 32844
rect 1162 32788 1230 32844
rect 1286 32788 1354 32844
rect 1410 32788 1478 32844
rect 1534 32788 1602 32844
rect 1658 32788 1726 32844
rect 1782 32788 1850 32844
rect 1906 32788 1916 32844
rect 104 32720 1916 32788
rect 104 32664 114 32720
rect 170 32664 238 32720
rect 294 32664 362 32720
rect 418 32664 486 32720
rect 542 32664 610 32720
rect 666 32664 734 32720
rect 790 32664 858 32720
rect 914 32664 982 32720
rect 1038 32664 1106 32720
rect 1162 32664 1230 32720
rect 1286 32664 1354 32720
rect 1410 32664 1478 32720
rect 1534 32664 1602 32720
rect 1658 32664 1726 32720
rect 1782 32664 1850 32720
rect 1906 32664 1916 32720
rect 104 32596 1916 32664
rect 104 32540 114 32596
rect 170 32540 238 32596
rect 294 32540 362 32596
rect 418 32540 486 32596
rect 542 32540 610 32596
rect 666 32540 734 32596
rect 790 32540 858 32596
rect 914 32540 982 32596
rect 1038 32540 1106 32596
rect 1162 32540 1230 32596
rect 1286 32540 1354 32596
rect 1410 32540 1478 32596
rect 1534 32540 1602 32596
rect 1658 32540 1726 32596
rect 1782 32540 1850 32596
rect 1906 32540 1916 32596
rect 104 32472 1916 32540
rect 104 32416 114 32472
rect 170 32416 238 32472
rect 294 32416 362 32472
rect 418 32416 486 32472
rect 542 32416 610 32472
rect 666 32416 734 32472
rect 790 32416 858 32472
rect 914 32416 982 32472
rect 1038 32416 1106 32472
rect 1162 32416 1230 32472
rect 1286 32416 1354 32472
rect 1410 32416 1478 32472
rect 1534 32416 1602 32472
rect 1658 32416 1726 32472
rect 1782 32416 1850 32472
rect 1906 32416 1916 32472
rect 104 32348 1916 32416
rect 104 32292 114 32348
rect 170 32292 238 32348
rect 294 32292 362 32348
rect 418 32292 486 32348
rect 542 32292 610 32348
rect 666 32292 734 32348
rect 790 32292 858 32348
rect 914 32292 982 32348
rect 1038 32292 1106 32348
rect 1162 32292 1230 32348
rect 1286 32292 1354 32348
rect 1410 32292 1478 32348
rect 1534 32292 1602 32348
rect 1658 32292 1726 32348
rect 1782 32292 1850 32348
rect 1906 32292 1916 32348
rect 104 32224 1916 32292
rect 104 32168 114 32224
rect 170 32168 238 32224
rect 294 32168 362 32224
rect 418 32168 486 32224
rect 542 32168 610 32224
rect 666 32168 734 32224
rect 790 32168 858 32224
rect 914 32168 982 32224
rect 1038 32168 1106 32224
rect 1162 32168 1230 32224
rect 1286 32168 1354 32224
rect 1410 32168 1478 32224
rect 1534 32168 1602 32224
rect 1658 32168 1726 32224
rect 1782 32168 1850 32224
rect 1906 32168 1916 32224
rect 104 32100 1916 32168
rect 104 32044 114 32100
rect 170 32044 238 32100
rect 294 32044 362 32100
rect 418 32044 486 32100
rect 542 32044 610 32100
rect 666 32044 734 32100
rect 790 32044 858 32100
rect 914 32044 982 32100
rect 1038 32044 1106 32100
rect 1162 32044 1230 32100
rect 1286 32044 1354 32100
rect 1410 32044 1478 32100
rect 1534 32044 1602 32100
rect 1658 32044 1726 32100
rect 1782 32044 1850 32100
rect 1906 32044 1916 32100
rect 104 31976 1916 32044
rect 104 31920 114 31976
rect 170 31920 238 31976
rect 294 31920 362 31976
rect 418 31920 486 31976
rect 542 31920 610 31976
rect 666 31920 734 31976
rect 790 31920 858 31976
rect 914 31920 982 31976
rect 1038 31920 1106 31976
rect 1162 31920 1230 31976
rect 1286 31920 1354 31976
rect 1410 31920 1478 31976
rect 1534 31920 1602 31976
rect 1658 31920 1726 31976
rect 1782 31920 1850 31976
rect 1906 31920 1916 31976
rect 104 31852 1916 31920
rect 104 31796 114 31852
rect 170 31796 238 31852
rect 294 31796 362 31852
rect 418 31796 486 31852
rect 542 31796 610 31852
rect 666 31796 734 31852
rect 790 31796 858 31852
rect 914 31796 982 31852
rect 1038 31796 1106 31852
rect 1162 31796 1230 31852
rect 1286 31796 1354 31852
rect 1410 31796 1478 31852
rect 1534 31796 1602 31852
rect 1658 31796 1726 31852
rect 1782 31796 1850 31852
rect 1906 31796 1916 31852
rect 104 31728 1916 31796
rect 104 31672 114 31728
rect 170 31672 238 31728
rect 294 31672 362 31728
rect 418 31672 486 31728
rect 542 31672 610 31728
rect 666 31672 734 31728
rect 790 31672 858 31728
rect 914 31672 982 31728
rect 1038 31672 1106 31728
rect 1162 31672 1230 31728
rect 1286 31672 1354 31728
rect 1410 31672 1478 31728
rect 1534 31672 1602 31728
rect 1658 31672 1726 31728
rect 1782 31672 1850 31728
rect 1906 31672 1916 31728
rect 104 31604 1916 31672
rect 104 31548 114 31604
rect 170 31548 238 31604
rect 294 31548 362 31604
rect 418 31548 486 31604
rect 542 31548 610 31604
rect 666 31548 734 31604
rect 790 31548 858 31604
rect 914 31548 982 31604
rect 1038 31548 1106 31604
rect 1162 31548 1230 31604
rect 1286 31548 1354 31604
rect 1410 31548 1478 31604
rect 1534 31548 1602 31604
rect 1658 31548 1726 31604
rect 1782 31548 1850 31604
rect 1906 31548 1916 31604
rect 104 31480 1916 31548
rect 104 31424 114 31480
rect 170 31424 238 31480
rect 294 31424 362 31480
rect 418 31424 486 31480
rect 542 31424 610 31480
rect 666 31424 734 31480
rect 790 31424 858 31480
rect 914 31424 982 31480
rect 1038 31424 1106 31480
rect 1162 31424 1230 31480
rect 1286 31424 1354 31480
rect 1410 31424 1478 31480
rect 1534 31424 1602 31480
rect 1658 31424 1726 31480
rect 1782 31424 1850 31480
rect 1906 31424 1916 31480
rect 104 31356 1916 31424
rect 104 31300 114 31356
rect 170 31300 238 31356
rect 294 31300 362 31356
rect 418 31300 486 31356
rect 542 31300 610 31356
rect 666 31300 734 31356
rect 790 31300 858 31356
rect 914 31300 982 31356
rect 1038 31300 1106 31356
rect 1162 31300 1230 31356
rect 1286 31300 1354 31356
rect 1410 31300 1478 31356
rect 1534 31300 1602 31356
rect 1658 31300 1726 31356
rect 1782 31300 1850 31356
rect 1906 31300 1916 31356
rect 104 31232 1916 31300
rect 104 31176 114 31232
rect 170 31176 238 31232
rect 294 31176 362 31232
rect 418 31176 486 31232
rect 542 31176 610 31232
rect 666 31176 734 31232
rect 790 31176 858 31232
rect 914 31176 982 31232
rect 1038 31176 1106 31232
rect 1162 31176 1230 31232
rect 1286 31176 1354 31232
rect 1410 31176 1478 31232
rect 1534 31176 1602 31232
rect 1658 31176 1726 31232
rect 1782 31176 1850 31232
rect 1906 31176 1916 31232
rect 104 31108 1916 31176
rect 104 31052 114 31108
rect 170 31052 238 31108
rect 294 31052 362 31108
rect 418 31052 486 31108
rect 542 31052 610 31108
rect 666 31052 734 31108
rect 790 31052 858 31108
rect 914 31052 982 31108
rect 1038 31052 1106 31108
rect 1162 31052 1230 31108
rect 1286 31052 1354 31108
rect 1410 31052 1478 31108
rect 1534 31052 1602 31108
rect 1658 31052 1726 31108
rect 1782 31052 1850 31108
rect 1906 31052 1916 31108
rect 104 30984 1916 31052
rect 104 30928 114 30984
rect 170 30928 238 30984
rect 294 30928 362 30984
rect 418 30928 486 30984
rect 542 30928 610 30984
rect 666 30928 734 30984
rect 790 30928 858 30984
rect 914 30928 982 30984
rect 1038 30928 1106 30984
rect 1162 30928 1230 30984
rect 1286 30928 1354 30984
rect 1410 30928 1478 30984
rect 1534 30928 1602 30984
rect 1658 30928 1726 30984
rect 1782 30928 1850 30984
rect 1906 30928 1916 30984
rect 104 30860 1916 30928
rect 104 30804 114 30860
rect 170 30804 238 30860
rect 294 30804 362 30860
rect 418 30804 486 30860
rect 542 30804 610 30860
rect 666 30804 734 30860
rect 790 30804 858 30860
rect 914 30804 982 30860
rect 1038 30804 1106 30860
rect 1162 30804 1230 30860
rect 1286 30804 1354 30860
rect 1410 30804 1478 30860
rect 1534 30804 1602 30860
rect 1658 30804 1726 30860
rect 1782 30804 1850 30860
rect 1906 30804 1916 30860
rect 104 30736 1916 30804
rect 104 30680 114 30736
rect 170 30680 238 30736
rect 294 30680 362 30736
rect 418 30680 486 30736
rect 542 30680 610 30736
rect 666 30680 734 30736
rect 790 30680 858 30736
rect 914 30680 982 30736
rect 1038 30680 1106 30736
rect 1162 30680 1230 30736
rect 1286 30680 1354 30736
rect 1410 30680 1478 30736
rect 1534 30680 1602 30736
rect 1658 30680 1726 30736
rect 1782 30680 1850 30736
rect 1906 30680 1916 30736
rect 104 30612 1916 30680
rect 104 30556 114 30612
rect 170 30556 238 30612
rect 294 30556 362 30612
rect 418 30556 486 30612
rect 542 30556 610 30612
rect 666 30556 734 30612
rect 790 30556 858 30612
rect 914 30556 982 30612
rect 1038 30556 1106 30612
rect 1162 30556 1230 30612
rect 1286 30556 1354 30612
rect 1410 30556 1478 30612
rect 1534 30556 1602 30612
rect 1658 30556 1726 30612
rect 1782 30556 1850 30612
rect 1906 30556 1916 30612
rect 104 30488 1916 30556
rect 104 30432 114 30488
rect 170 30432 238 30488
rect 294 30432 362 30488
rect 418 30432 486 30488
rect 542 30432 610 30488
rect 666 30432 734 30488
rect 790 30432 858 30488
rect 914 30432 982 30488
rect 1038 30432 1106 30488
rect 1162 30432 1230 30488
rect 1286 30432 1354 30488
rect 1410 30432 1478 30488
rect 1534 30432 1602 30488
rect 1658 30432 1726 30488
rect 1782 30432 1850 30488
rect 1906 30432 1916 30488
rect 104 30364 1916 30432
rect 104 30308 114 30364
rect 170 30308 238 30364
rect 294 30308 362 30364
rect 418 30308 486 30364
rect 542 30308 610 30364
rect 666 30308 734 30364
rect 790 30308 858 30364
rect 914 30308 982 30364
rect 1038 30308 1106 30364
rect 1162 30308 1230 30364
rect 1286 30308 1354 30364
rect 1410 30308 1478 30364
rect 1534 30308 1602 30364
rect 1658 30308 1726 30364
rect 1782 30308 1850 30364
rect 1906 30308 1916 30364
rect 104 30240 1916 30308
rect 104 30184 114 30240
rect 170 30184 238 30240
rect 294 30184 362 30240
rect 418 30184 486 30240
rect 542 30184 610 30240
rect 666 30184 734 30240
rect 790 30184 858 30240
rect 914 30184 982 30240
rect 1038 30184 1106 30240
rect 1162 30184 1230 30240
rect 1286 30184 1354 30240
rect 1410 30184 1478 30240
rect 1534 30184 1602 30240
rect 1658 30184 1726 30240
rect 1782 30184 1850 30240
rect 1906 30184 1916 30240
rect 104 30174 1916 30184
rect 104 29643 1916 29653
rect 104 29587 114 29643
rect 170 29587 238 29643
rect 294 29587 362 29643
rect 418 29587 486 29643
rect 542 29587 610 29643
rect 666 29587 734 29643
rect 790 29587 858 29643
rect 914 29587 982 29643
rect 1038 29587 1106 29643
rect 1162 29587 1230 29643
rect 1286 29587 1354 29643
rect 1410 29587 1478 29643
rect 1534 29587 1602 29643
rect 1658 29587 1726 29643
rect 1782 29587 1850 29643
rect 1906 29587 1916 29643
rect 104 29519 1916 29587
rect 104 29463 114 29519
rect 170 29463 238 29519
rect 294 29463 362 29519
rect 418 29463 486 29519
rect 542 29463 610 29519
rect 666 29463 734 29519
rect 790 29463 858 29519
rect 914 29463 982 29519
rect 1038 29463 1106 29519
rect 1162 29463 1230 29519
rect 1286 29463 1354 29519
rect 1410 29463 1478 29519
rect 1534 29463 1602 29519
rect 1658 29463 1726 29519
rect 1782 29463 1850 29519
rect 1906 29463 1916 29519
rect 104 29395 1916 29463
rect 104 29339 114 29395
rect 170 29339 238 29395
rect 294 29339 362 29395
rect 418 29339 486 29395
rect 542 29339 610 29395
rect 666 29339 734 29395
rect 790 29339 858 29395
rect 914 29339 982 29395
rect 1038 29339 1106 29395
rect 1162 29339 1230 29395
rect 1286 29339 1354 29395
rect 1410 29339 1478 29395
rect 1534 29339 1602 29395
rect 1658 29339 1726 29395
rect 1782 29339 1850 29395
rect 1906 29339 1916 29395
rect 104 29271 1916 29339
rect 104 29215 114 29271
rect 170 29215 238 29271
rect 294 29215 362 29271
rect 418 29215 486 29271
rect 542 29215 610 29271
rect 666 29215 734 29271
rect 790 29215 858 29271
rect 914 29215 982 29271
rect 1038 29215 1106 29271
rect 1162 29215 1230 29271
rect 1286 29215 1354 29271
rect 1410 29215 1478 29271
rect 1534 29215 1602 29271
rect 1658 29215 1726 29271
rect 1782 29215 1850 29271
rect 1906 29215 1916 29271
rect 104 29147 1916 29215
rect 104 29091 114 29147
rect 170 29091 238 29147
rect 294 29091 362 29147
rect 418 29091 486 29147
rect 542 29091 610 29147
rect 666 29091 734 29147
rect 790 29091 858 29147
rect 914 29091 982 29147
rect 1038 29091 1106 29147
rect 1162 29091 1230 29147
rect 1286 29091 1354 29147
rect 1410 29091 1478 29147
rect 1534 29091 1602 29147
rect 1658 29091 1726 29147
rect 1782 29091 1850 29147
rect 1906 29091 1916 29147
rect 104 29023 1916 29091
rect 104 28967 114 29023
rect 170 28967 238 29023
rect 294 28967 362 29023
rect 418 28967 486 29023
rect 542 28967 610 29023
rect 666 28967 734 29023
rect 790 28967 858 29023
rect 914 28967 982 29023
rect 1038 28967 1106 29023
rect 1162 28967 1230 29023
rect 1286 28967 1354 29023
rect 1410 28967 1478 29023
rect 1534 28967 1602 29023
rect 1658 28967 1726 29023
rect 1782 28967 1850 29023
rect 1906 28967 1916 29023
rect 104 28899 1916 28967
rect 104 28843 114 28899
rect 170 28843 238 28899
rect 294 28843 362 28899
rect 418 28843 486 28899
rect 542 28843 610 28899
rect 666 28843 734 28899
rect 790 28843 858 28899
rect 914 28843 982 28899
rect 1038 28843 1106 28899
rect 1162 28843 1230 28899
rect 1286 28843 1354 28899
rect 1410 28843 1478 28899
rect 1534 28843 1602 28899
rect 1658 28843 1726 28899
rect 1782 28843 1850 28899
rect 1906 28843 1916 28899
rect 104 28775 1916 28843
rect 104 28719 114 28775
rect 170 28719 238 28775
rect 294 28719 362 28775
rect 418 28719 486 28775
rect 542 28719 610 28775
rect 666 28719 734 28775
rect 790 28719 858 28775
rect 914 28719 982 28775
rect 1038 28719 1106 28775
rect 1162 28719 1230 28775
rect 1286 28719 1354 28775
rect 1410 28719 1478 28775
rect 1534 28719 1602 28775
rect 1658 28719 1726 28775
rect 1782 28719 1850 28775
rect 1906 28719 1916 28775
rect 104 28651 1916 28719
rect 104 28595 114 28651
rect 170 28595 238 28651
rect 294 28595 362 28651
rect 418 28595 486 28651
rect 542 28595 610 28651
rect 666 28595 734 28651
rect 790 28595 858 28651
rect 914 28595 982 28651
rect 1038 28595 1106 28651
rect 1162 28595 1230 28651
rect 1286 28595 1354 28651
rect 1410 28595 1478 28651
rect 1534 28595 1602 28651
rect 1658 28595 1726 28651
rect 1782 28595 1850 28651
rect 1906 28595 1916 28651
rect 104 28527 1916 28595
rect 104 28471 114 28527
rect 170 28471 238 28527
rect 294 28471 362 28527
rect 418 28471 486 28527
rect 542 28471 610 28527
rect 666 28471 734 28527
rect 790 28471 858 28527
rect 914 28471 982 28527
rect 1038 28471 1106 28527
rect 1162 28471 1230 28527
rect 1286 28471 1354 28527
rect 1410 28471 1478 28527
rect 1534 28471 1602 28527
rect 1658 28471 1726 28527
rect 1782 28471 1850 28527
rect 1906 28471 1916 28527
rect 104 28403 1916 28471
rect 104 28347 114 28403
rect 170 28347 238 28403
rect 294 28347 362 28403
rect 418 28347 486 28403
rect 542 28347 610 28403
rect 666 28347 734 28403
rect 790 28347 858 28403
rect 914 28347 982 28403
rect 1038 28347 1106 28403
rect 1162 28347 1230 28403
rect 1286 28347 1354 28403
rect 1410 28347 1478 28403
rect 1534 28347 1602 28403
rect 1658 28347 1726 28403
rect 1782 28347 1850 28403
rect 1906 28347 1916 28403
rect 104 28279 1916 28347
rect 104 28223 114 28279
rect 170 28223 238 28279
rect 294 28223 362 28279
rect 418 28223 486 28279
rect 542 28223 610 28279
rect 666 28223 734 28279
rect 790 28223 858 28279
rect 914 28223 982 28279
rect 1038 28223 1106 28279
rect 1162 28223 1230 28279
rect 1286 28223 1354 28279
rect 1410 28223 1478 28279
rect 1534 28223 1602 28279
rect 1658 28223 1726 28279
rect 1782 28223 1850 28279
rect 1906 28223 1916 28279
rect 104 28155 1916 28223
rect 104 28099 114 28155
rect 170 28099 238 28155
rect 294 28099 362 28155
rect 418 28099 486 28155
rect 542 28099 610 28155
rect 666 28099 734 28155
rect 790 28099 858 28155
rect 914 28099 982 28155
rect 1038 28099 1106 28155
rect 1162 28099 1230 28155
rect 1286 28099 1354 28155
rect 1410 28099 1478 28155
rect 1534 28099 1602 28155
rect 1658 28099 1726 28155
rect 1782 28099 1850 28155
rect 1906 28099 1916 28155
rect 104 28031 1916 28099
rect 104 27975 114 28031
rect 170 27975 238 28031
rect 294 27975 362 28031
rect 418 27975 486 28031
rect 542 27975 610 28031
rect 666 27975 734 28031
rect 790 27975 858 28031
rect 914 27975 982 28031
rect 1038 27975 1106 28031
rect 1162 27975 1230 28031
rect 1286 27975 1354 28031
rect 1410 27975 1478 28031
rect 1534 27975 1602 28031
rect 1658 27975 1726 28031
rect 1782 27975 1850 28031
rect 1906 27975 1916 28031
rect 104 27907 1916 27975
rect 104 27851 114 27907
rect 170 27851 238 27907
rect 294 27851 362 27907
rect 418 27851 486 27907
rect 542 27851 610 27907
rect 666 27851 734 27907
rect 790 27851 858 27907
rect 914 27851 982 27907
rect 1038 27851 1106 27907
rect 1162 27851 1230 27907
rect 1286 27851 1354 27907
rect 1410 27851 1478 27907
rect 1534 27851 1602 27907
rect 1658 27851 1726 27907
rect 1782 27851 1850 27907
rect 1906 27851 1916 27907
rect 104 27783 1916 27851
rect 104 27727 114 27783
rect 170 27727 238 27783
rect 294 27727 362 27783
rect 418 27727 486 27783
rect 542 27727 610 27783
rect 666 27727 734 27783
rect 790 27727 858 27783
rect 914 27727 982 27783
rect 1038 27727 1106 27783
rect 1162 27727 1230 27783
rect 1286 27727 1354 27783
rect 1410 27727 1478 27783
rect 1534 27727 1602 27783
rect 1658 27727 1726 27783
rect 1782 27727 1850 27783
rect 1906 27727 1916 27783
rect 104 27659 1916 27727
rect 104 27603 114 27659
rect 170 27603 238 27659
rect 294 27603 362 27659
rect 418 27603 486 27659
rect 542 27603 610 27659
rect 666 27603 734 27659
rect 790 27603 858 27659
rect 914 27603 982 27659
rect 1038 27603 1106 27659
rect 1162 27603 1230 27659
rect 1286 27603 1354 27659
rect 1410 27603 1478 27659
rect 1534 27603 1602 27659
rect 1658 27603 1726 27659
rect 1782 27603 1850 27659
rect 1906 27603 1916 27659
rect 104 27535 1916 27603
rect 104 27479 114 27535
rect 170 27479 238 27535
rect 294 27479 362 27535
rect 418 27479 486 27535
rect 542 27479 610 27535
rect 666 27479 734 27535
rect 790 27479 858 27535
rect 914 27479 982 27535
rect 1038 27479 1106 27535
rect 1162 27479 1230 27535
rect 1286 27479 1354 27535
rect 1410 27479 1478 27535
rect 1534 27479 1602 27535
rect 1658 27479 1726 27535
rect 1782 27479 1850 27535
rect 1906 27479 1916 27535
rect 104 27411 1916 27479
rect 104 27355 114 27411
rect 170 27355 238 27411
rect 294 27355 362 27411
rect 418 27355 486 27411
rect 542 27355 610 27411
rect 666 27355 734 27411
rect 790 27355 858 27411
rect 914 27355 982 27411
rect 1038 27355 1106 27411
rect 1162 27355 1230 27411
rect 1286 27355 1354 27411
rect 1410 27355 1478 27411
rect 1534 27355 1602 27411
rect 1658 27355 1726 27411
rect 1782 27355 1850 27411
rect 1906 27355 1916 27411
rect 104 27287 1916 27355
rect 104 27231 114 27287
rect 170 27231 238 27287
rect 294 27231 362 27287
rect 418 27231 486 27287
rect 542 27231 610 27287
rect 666 27231 734 27287
rect 790 27231 858 27287
rect 914 27231 982 27287
rect 1038 27231 1106 27287
rect 1162 27231 1230 27287
rect 1286 27231 1354 27287
rect 1410 27231 1478 27287
rect 1534 27231 1602 27287
rect 1658 27231 1726 27287
rect 1782 27231 1850 27287
rect 1906 27231 1916 27287
rect 104 27163 1916 27231
rect 104 27107 114 27163
rect 170 27107 238 27163
rect 294 27107 362 27163
rect 418 27107 486 27163
rect 542 27107 610 27163
rect 666 27107 734 27163
rect 790 27107 858 27163
rect 914 27107 982 27163
rect 1038 27107 1106 27163
rect 1162 27107 1230 27163
rect 1286 27107 1354 27163
rect 1410 27107 1478 27163
rect 1534 27107 1602 27163
rect 1658 27107 1726 27163
rect 1782 27107 1850 27163
rect 1906 27107 1916 27163
rect 104 27039 1916 27107
rect 104 26983 114 27039
rect 170 26983 238 27039
rect 294 26983 362 27039
rect 418 26983 486 27039
rect 542 26983 610 27039
rect 666 26983 734 27039
rect 790 26983 858 27039
rect 914 26983 982 27039
rect 1038 26983 1106 27039
rect 1162 26983 1230 27039
rect 1286 26983 1354 27039
rect 1410 26983 1478 27039
rect 1534 26983 1602 27039
rect 1658 26983 1726 27039
rect 1782 26983 1850 27039
rect 1906 26983 1916 27039
rect 104 26973 1916 26983
rect 104 26501 1916 26511
rect 104 26445 114 26501
rect 170 26445 238 26501
rect 294 26445 362 26501
rect 418 26445 486 26501
rect 542 26445 610 26501
rect 666 26445 734 26501
rect 790 26445 858 26501
rect 914 26445 982 26501
rect 1038 26445 1106 26501
rect 1162 26445 1230 26501
rect 1286 26445 1354 26501
rect 1410 26445 1478 26501
rect 1534 26445 1602 26501
rect 1658 26445 1726 26501
rect 1782 26445 1850 26501
rect 1906 26445 1916 26501
rect 104 26377 1916 26445
rect 104 26321 114 26377
rect 170 26321 238 26377
rect 294 26321 362 26377
rect 418 26321 486 26377
rect 542 26321 610 26377
rect 666 26321 734 26377
rect 790 26321 858 26377
rect 914 26321 982 26377
rect 1038 26321 1106 26377
rect 1162 26321 1230 26377
rect 1286 26321 1354 26377
rect 1410 26321 1478 26377
rect 1534 26321 1602 26377
rect 1658 26321 1726 26377
rect 1782 26321 1850 26377
rect 1906 26321 1916 26377
rect 104 26253 1916 26321
rect 104 26197 114 26253
rect 170 26197 238 26253
rect 294 26197 362 26253
rect 418 26197 486 26253
rect 542 26197 610 26253
rect 666 26197 734 26253
rect 790 26197 858 26253
rect 914 26197 982 26253
rect 1038 26197 1106 26253
rect 1162 26197 1230 26253
rect 1286 26197 1354 26253
rect 1410 26197 1478 26253
rect 1534 26197 1602 26253
rect 1658 26197 1726 26253
rect 1782 26197 1850 26253
rect 1906 26197 1916 26253
rect 104 26129 1916 26197
rect 104 26073 114 26129
rect 170 26073 238 26129
rect 294 26073 362 26129
rect 418 26073 486 26129
rect 542 26073 610 26129
rect 666 26073 734 26129
rect 790 26073 858 26129
rect 914 26073 982 26129
rect 1038 26073 1106 26129
rect 1162 26073 1230 26129
rect 1286 26073 1354 26129
rect 1410 26073 1478 26129
rect 1534 26073 1602 26129
rect 1658 26073 1726 26129
rect 1782 26073 1850 26129
rect 1906 26073 1916 26129
rect 104 26005 1916 26073
rect 104 25949 114 26005
rect 170 25949 238 26005
rect 294 25949 362 26005
rect 418 25949 486 26005
rect 542 25949 610 26005
rect 666 25949 734 26005
rect 790 25949 858 26005
rect 914 25949 982 26005
rect 1038 25949 1106 26005
rect 1162 25949 1230 26005
rect 1286 25949 1354 26005
rect 1410 25949 1478 26005
rect 1534 25949 1602 26005
rect 1658 25949 1726 26005
rect 1782 25949 1850 26005
rect 1906 25949 1916 26005
rect 104 25881 1916 25949
rect 104 25825 114 25881
rect 170 25825 238 25881
rect 294 25825 362 25881
rect 418 25825 486 25881
rect 542 25825 610 25881
rect 666 25825 734 25881
rect 790 25825 858 25881
rect 914 25825 982 25881
rect 1038 25825 1106 25881
rect 1162 25825 1230 25881
rect 1286 25825 1354 25881
rect 1410 25825 1478 25881
rect 1534 25825 1602 25881
rect 1658 25825 1726 25881
rect 1782 25825 1850 25881
rect 1906 25825 1916 25881
rect 104 25757 1916 25825
rect 104 25701 114 25757
rect 170 25701 238 25757
rect 294 25701 362 25757
rect 418 25701 486 25757
rect 542 25701 610 25757
rect 666 25701 734 25757
rect 790 25701 858 25757
rect 914 25701 982 25757
rect 1038 25701 1106 25757
rect 1162 25701 1230 25757
rect 1286 25701 1354 25757
rect 1410 25701 1478 25757
rect 1534 25701 1602 25757
rect 1658 25701 1726 25757
rect 1782 25701 1850 25757
rect 1906 25701 1916 25757
rect 104 25633 1916 25701
rect 104 25577 114 25633
rect 170 25577 238 25633
rect 294 25577 362 25633
rect 418 25577 486 25633
rect 542 25577 610 25633
rect 666 25577 734 25633
rect 790 25577 858 25633
rect 914 25577 982 25633
rect 1038 25577 1106 25633
rect 1162 25577 1230 25633
rect 1286 25577 1354 25633
rect 1410 25577 1478 25633
rect 1534 25577 1602 25633
rect 1658 25577 1726 25633
rect 1782 25577 1850 25633
rect 1906 25577 1916 25633
rect 104 25509 1916 25577
rect 104 25453 114 25509
rect 170 25453 238 25509
rect 294 25453 362 25509
rect 418 25453 486 25509
rect 542 25453 610 25509
rect 666 25453 734 25509
rect 790 25453 858 25509
rect 914 25453 982 25509
rect 1038 25453 1106 25509
rect 1162 25453 1230 25509
rect 1286 25453 1354 25509
rect 1410 25453 1478 25509
rect 1534 25453 1602 25509
rect 1658 25453 1726 25509
rect 1782 25453 1850 25509
rect 1906 25453 1916 25509
rect 104 25385 1916 25453
rect 104 25329 114 25385
rect 170 25329 238 25385
rect 294 25329 362 25385
rect 418 25329 486 25385
rect 542 25329 610 25385
rect 666 25329 734 25385
rect 790 25329 858 25385
rect 914 25329 982 25385
rect 1038 25329 1106 25385
rect 1162 25329 1230 25385
rect 1286 25329 1354 25385
rect 1410 25329 1478 25385
rect 1534 25329 1602 25385
rect 1658 25329 1726 25385
rect 1782 25329 1850 25385
rect 1906 25329 1916 25385
rect 104 25319 1916 25329
rect 104 24888 1916 24898
rect 104 24832 114 24888
rect 170 24832 238 24888
rect 294 24832 362 24888
rect 418 24832 486 24888
rect 542 24832 610 24888
rect 666 24832 734 24888
rect 790 24832 858 24888
rect 914 24832 982 24888
rect 1038 24832 1106 24888
rect 1162 24832 1230 24888
rect 1286 24832 1354 24888
rect 1410 24832 1478 24888
rect 1534 24832 1602 24888
rect 1658 24832 1726 24888
rect 1782 24832 1850 24888
rect 1906 24832 1916 24888
rect 104 24764 1916 24832
rect 104 24708 114 24764
rect 170 24708 238 24764
rect 294 24708 362 24764
rect 418 24708 486 24764
rect 542 24708 610 24764
rect 666 24708 734 24764
rect 790 24708 858 24764
rect 914 24708 982 24764
rect 1038 24708 1106 24764
rect 1162 24708 1230 24764
rect 1286 24708 1354 24764
rect 1410 24708 1478 24764
rect 1534 24708 1602 24764
rect 1658 24708 1726 24764
rect 1782 24708 1850 24764
rect 1906 24708 1916 24764
rect 104 24640 1916 24708
rect 104 24584 114 24640
rect 170 24584 238 24640
rect 294 24584 362 24640
rect 418 24584 486 24640
rect 542 24584 610 24640
rect 666 24584 734 24640
rect 790 24584 858 24640
rect 914 24584 982 24640
rect 1038 24584 1106 24640
rect 1162 24584 1230 24640
rect 1286 24584 1354 24640
rect 1410 24584 1478 24640
rect 1534 24584 1602 24640
rect 1658 24584 1726 24640
rect 1782 24584 1850 24640
rect 1906 24584 1916 24640
rect 104 24516 1916 24584
rect 104 24460 114 24516
rect 170 24460 238 24516
rect 294 24460 362 24516
rect 418 24460 486 24516
rect 542 24460 610 24516
rect 666 24460 734 24516
rect 790 24460 858 24516
rect 914 24460 982 24516
rect 1038 24460 1106 24516
rect 1162 24460 1230 24516
rect 1286 24460 1354 24516
rect 1410 24460 1478 24516
rect 1534 24460 1602 24516
rect 1658 24460 1726 24516
rect 1782 24460 1850 24516
rect 1906 24460 1916 24516
rect 104 24392 1916 24460
rect 104 24336 114 24392
rect 170 24336 238 24392
rect 294 24336 362 24392
rect 418 24336 486 24392
rect 542 24336 610 24392
rect 666 24336 734 24392
rect 790 24336 858 24392
rect 914 24336 982 24392
rect 1038 24336 1106 24392
rect 1162 24336 1230 24392
rect 1286 24336 1354 24392
rect 1410 24336 1478 24392
rect 1534 24336 1602 24392
rect 1658 24336 1726 24392
rect 1782 24336 1850 24392
rect 1906 24336 1916 24392
rect 104 24268 1916 24336
rect 104 24212 114 24268
rect 170 24212 238 24268
rect 294 24212 362 24268
rect 418 24212 486 24268
rect 542 24212 610 24268
rect 666 24212 734 24268
rect 790 24212 858 24268
rect 914 24212 982 24268
rect 1038 24212 1106 24268
rect 1162 24212 1230 24268
rect 1286 24212 1354 24268
rect 1410 24212 1478 24268
rect 1534 24212 1602 24268
rect 1658 24212 1726 24268
rect 1782 24212 1850 24268
rect 1906 24212 1916 24268
rect 104 24144 1916 24212
rect 104 24088 114 24144
rect 170 24088 238 24144
rect 294 24088 362 24144
rect 418 24088 486 24144
rect 542 24088 610 24144
rect 666 24088 734 24144
rect 790 24088 858 24144
rect 914 24088 982 24144
rect 1038 24088 1106 24144
rect 1162 24088 1230 24144
rect 1286 24088 1354 24144
rect 1410 24088 1478 24144
rect 1534 24088 1602 24144
rect 1658 24088 1726 24144
rect 1782 24088 1850 24144
rect 1906 24088 1916 24144
rect 104 24020 1916 24088
rect 104 23964 114 24020
rect 170 23964 238 24020
rect 294 23964 362 24020
rect 418 23964 486 24020
rect 542 23964 610 24020
rect 666 23964 734 24020
rect 790 23964 858 24020
rect 914 23964 982 24020
rect 1038 23964 1106 24020
rect 1162 23964 1230 24020
rect 1286 23964 1354 24020
rect 1410 23964 1478 24020
rect 1534 23964 1602 24020
rect 1658 23964 1726 24020
rect 1782 23964 1850 24020
rect 1906 23964 1916 24020
rect 104 23896 1916 23964
rect 104 23840 114 23896
rect 170 23840 238 23896
rect 294 23840 362 23896
rect 418 23840 486 23896
rect 542 23840 610 23896
rect 666 23840 734 23896
rect 790 23840 858 23896
rect 914 23840 982 23896
rect 1038 23840 1106 23896
rect 1162 23840 1230 23896
rect 1286 23840 1354 23896
rect 1410 23840 1478 23896
rect 1534 23840 1602 23896
rect 1658 23840 1726 23896
rect 1782 23840 1850 23896
rect 1906 23840 1916 23896
rect 104 23772 1916 23840
rect 104 23716 114 23772
rect 170 23716 238 23772
rect 294 23716 362 23772
rect 418 23716 486 23772
rect 542 23716 610 23772
rect 666 23716 734 23772
rect 790 23716 858 23772
rect 914 23716 982 23772
rect 1038 23716 1106 23772
rect 1162 23716 1230 23772
rect 1286 23716 1354 23772
rect 1410 23716 1478 23772
rect 1534 23716 1602 23772
rect 1658 23716 1726 23772
rect 1782 23716 1850 23772
rect 1906 23716 1916 23772
rect 104 23706 1916 23716
rect 104 23234 1916 23244
rect 104 23178 114 23234
rect 170 23178 238 23234
rect 294 23178 362 23234
rect 418 23178 486 23234
rect 542 23178 610 23234
rect 666 23178 734 23234
rect 790 23178 858 23234
rect 914 23178 982 23234
rect 1038 23178 1106 23234
rect 1162 23178 1230 23234
rect 1286 23178 1354 23234
rect 1410 23178 1478 23234
rect 1534 23178 1602 23234
rect 1658 23178 1726 23234
rect 1782 23178 1850 23234
rect 1906 23178 1916 23234
rect 104 23110 1916 23178
rect 104 23054 114 23110
rect 170 23054 238 23110
rect 294 23054 362 23110
rect 418 23054 486 23110
rect 542 23054 610 23110
rect 666 23054 734 23110
rect 790 23054 858 23110
rect 914 23054 982 23110
rect 1038 23054 1106 23110
rect 1162 23054 1230 23110
rect 1286 23054 1354 23110
rect 1410 23054 1478 23110
rect 1534 23054 1602 23110
rect 1658 23054 1726 23110
rect 1782 23054 1850 23110
rect 1906 23054 1916 23110
rect 104 22986 1916 23054
rect 104 22930 114 22986
rect 170 22930 238 22986
rect 294 22930 362 22986
rect 418 22930 486 22986
rect 542 22930 610 22986
rect 666 22930 734 22986
rect 790 22930 858 22986
rect 914 22930 982 22986
rect 1038 22930 1106 22986
rect 1162 22930 1230 22986
rect 1286 22930 1354 22986
rect 1410 22930 1478 22986
rect 1534 22930 1602 22986
rect 1658 22930 1726 22986
rect 1782 22930 1850 22986
rect 1906 22930 1916 22986
rect 104 22862 1916 22930
rect 104 22806 114 22862
rect 170 22806 238 22862
rect 294 22806 362 22862
rect 418 22806 486 22862
rect 542 22806 610 22862
rect 666 22806 734 22862
rect 790 22806 858 22862
rect 914 22806 982 22862
rect 1038 22806 1106 22862
rect 1162 22806 1230 22862
rect 1286 22806 1354 22862
rect 1410 22806 1478 22862
rect 1534 22806 1602 22862
rect 1658 22806 1726 22862
rect 1782 22806 1850 22862
rect 1906 22806 1916 22862
rect 104 22738 1916 22806
rect 104 22682 114 22738
rect 170 22682 238 22738
rect 294 22682 362 22738
rect 418 22682 486 22738
rect 542 22682 610 22738
rect 666 22682 734 22738
rect 790 22682 858 22738
rect 914 22682 982 22738
rect 1038 22682 1106 22738
rect 1162 22682 1230 22738
rect 1286 22682 1354 22738
rect 1410 22682 1478 22738
rect 1534 22682 1602 22738
rect 1658 22682 1726 22738
rect 1782 22682 1850 22738
rect 1906 22682 1916 22738
rect 104 22614 1916 22682
rect 104 22558 114 22614
rect 170 22558 238 22614
rect 294 22558 362 22614
rect 418 22558 486 22614
rect 542 22558 610 22614
rect 666 22558 734 22614
rect 790 22558 858 22614
rect 914 22558 982 22614
rect 1038 22558 1106 22614
rect 1162 22558 1230 22614
rect 1286 22558 1354 22614
rect 1410 22558 1478 22614
rect 1534 22558 1602 22614
rect 1658 22558 1726 22614
rect 1782 22558 1850 22614
rect 1906 22558 1916 22614
rect 104 22490 1916 22558
rect 104 22434 114 22490
rect 170 22434 238 22490
rect 294 22434 362 22490
rect 418 22434 486 22490
rect 542 22434 610 22490
rect 666 22434 734 22490
rect 790 22434 858 22490
rect 914 22434 982 22490
rect 1038 22434 1106 22490
rect 1162 22434 1230 22490
rect 1286 22434 1354 22490
rect 1410 22434 1478 22490
rect 1534 22434 1602 22490
rect 1658 22434 1726 22490
rect 1782 22434 1850 22490
rect 1906 22434 1916 22490
rect 104 22366 1916 22434
rect 104 22310 114 22366
rect 170 22310 238 22366
rect 294 22310 362 22366
rect 418 22310 486 22366
rect 542 22310 610 22366
rect 666 22310 734 22366
rect 790 22310 858 22366
rect 914 22310 982 22366
rect 1038 22310 1106 22366
rect 1162 22310 1230 22366
rect 1286 22310 1354 22366
rect 1410 22310 1478 22366
rect 1534 22310 1602 22366
rect 1658 22310 1726 22366
rect 1782 22310 1850 22366
rect 1906 22310 1916 22366
rect 104 22242 1916 22310
rect 104 22186 114 22242
rect 170 22186 238 22242
rect 294 22186 362 22242
rect 418 22186 486 22242
rect 542 22186 610 22242
rect 666 22186 734 22242
rect 790 22186 858 22242
rect 914 22186 982 22242
rect 1038 22186 1106 22242
rect 1162 22186 1230 22242
rect 1286 22186 1354 22242
rect 1410 22186 1478 22242
rect 1534 22186 1602 22242
rect 1658 22186 1726 22242
rect 1782 22186 1850 22242
rect 1906 22186 1916 22242
rect 104 22118 1916 22186
rect 104 22062 114 22118
rect 170 22062 238 22118
rect 294 22062 362 22118
rect 418 22062 486 22118
rect 542 22062 610 22118
rect 666 22062 734 22118
rect 790 22062 858 22118
rect 914 22062 982 22118
rect 1038 22062 1106 22118
rect 1162 22062 1230 22118
rect 1286 22062 1354 22118
rect 1410 22062 1478 22118
rect 1534 22062 1602 22118
rect 1658 22062 1726 22118
rect 1782 22062 1850 22118
rect 1906 22062 1916 22118
rect 104 21994 1916 22062
rect 104 21938 114 21994
rect 170 21938 238 21994
rect 294 21938 362 21994
rect 418 21938 486 21994
rect 542 21938 610 21994
rect 666 21938 734 21994
rect 790 21938 858 21994
rect 914 21938 982 21994
rect 1038 21938 1106 21994
rect 1162 21938 1230 21994
rect 1286 21938 1354 21994
rect 1410 21938 1478 21994
rect 1534 21938 1602 21994
rect 1658 21938 1726 21994
rect 1782 21938 1850 21994
rect 1906 21938 1916 21994
rect 104 21870 1916 21938
rect 104 21814 114 21870
rect 170 21814 238 21870
rect 294 21814 362 21870
rect 418 21814 486 21870
rect 542 21814 610 21870
rect 666 21814 734 21870
rect 790 21814 858 21870
rect 914 21814 982 21870
rect 1038 21814 1106 21870
rect 1162 21814 1230 21870
rect 1286 21814 1354 21870
rect 1410 21814 1478 21870
rect 1534 21814 1602 21870
rect 1658 21814 1726 21870
rect 1782 21814 1850 21870
rect 1906 21814 1916 21870
rect 104 21746 1916 21814
rect 104 21690 114 21746
rect 170 21690 238 21746
rect 294 21690 362 21746
rect 418 21690 486 21746
rect 542 21690 610 21746
rect 666 21690 734 21746
rect 790 21690 858 21746
rect 914 21690 982 21746
rect 1038 21690 1106 21746
rect 1162 21690 1230 21746
rect 1286 21690 1354 21746
rect 1410 21690 1478 21746
rect 1534 21690 1602 21746
rect 1658 21690 1726 21746
rect 1782 21690 1850 21746
rect 1906 21690 1916 21746
rect 104 21622 1916 21690
rect 104 21566 114 21622
rect 170 21566 238 21622
rect 294 21566 362 21622
rect 418 21566 486 21622
rect 542 21566 610 21622
rect 666 21566 734 21622
rect 790 21566 858 21622
rect 914 21566 982 21622
rect 1038 21566 1106 21622
rect 1162 21566 1230 21622
rect 1286 21566 1354 21622
rect 1410 21566 1478 21622
rect 1534 21566 1602 21622
rect 1658 21566 1726 21622
rect 1782 21566 1850 21622
rect 1906 21566 1916 21622
rect 104 21498 1916 21566
rect 104 21442 114 21498
rect 170 21442 238 21498
rect 294 21442 362 21498
rect 418 21442 486 21498
rect 542 21442 610 21498
rect 666 21442 734 21498
rect 790 21442 858 21498
rect 914 21442 982 21498
rect 1038 21442 1106 21498
rect 1162 21442 1230 21498
rect 1286 21442 1354 21498
rect 1410 21442 1478 21498
rect 1534 21442 1602 21498
rect 1658 21442 1726 21498
rect 1782 21442 1850 21498
rect 1906 21442 1916 21498
rect 104 21374 1916 21442
rect 104 21318 114 21374
rect 170 21318 238 21374
rect 294 21318 362 21374
rect 418 21318 486 21374
rect 542 21318 610 21374
rect 666 21318 734 21374
rect 790 21318 858 21374
rect 914 21318 982 21374
rect 1038 21318 1106 21374
rect 1162 21318 1230 21374
rect 1286 21318 1354 21374
rect 1410 21318 1478 21374
rect 1534 21318 1602 21374
rect 1658 21318 1726 21374
rect 1782 21318 1850 21374
rect 1906 21318 1916 21374
rect 104 21250 1916 21318
rect 104 21194 114 21250
rect 170 21194 238 21250
rect 294 21194 362 21250
rect 418 21194 486 21250
rect 542 21194 610 21250
rect 666 21194 734 21250
rect 790 21194 858 21250
rect 914 21194 982 21250
rect 1038 21194 1106 21250
rect 1162 21194 1230 21250
rect 1286 21194 1354 21250
rect 1410 21194 1478 21250
rect 1534 21194 1602 21250
rect 1658 21194 1726 21250
rect 1782 21194 1850 21250
rect 1906 21194 1916 21250
rect 104 21126 1916 21194
rect 104 21070 114 21126
rect 170 21070 238 21126
rect 294 21070 362 21126
rect 418 21070 486 21126
rect 542 21070 610 21126
rect 666 21070 734 21126
rect 790 21070 858 21126
rect 914 21070 982 21126
rect 1038 21070 1106 21126
rect 1162 21070 1230 21126
rect 1286 21070 1354 21126
rect 1410 21070 1478 21126
rect 1534 21070 1602 21126
rect 1658 21070 1726 21126
rect 1782 21070 1850 21126
rect 1906 21070 1916 21126
rect 104 21002 1916 21070
rect 104 20946 114 21002
rect 170 20946 238 21002
rect 294 20946 362 21002
rect 418 20946 486 21002
rect 542 20946 610 21002
rect 666 20946 734 21002
rect 790 20946 858 21002
rect 914 20946 982 21002
rect 1038 20946 1106 21002
rect 1162 20946 1230 21002
rect 1286 20946 1354 21002
rect 1410 20946 1478 21002
rect 1534 20946 1602 21002
rect 1658 20946 1726 21002
rect 1782 20946 1850 21002
rect 1906 20946 1916 21002
rect 104 20878 1916 20946
rect 104 20822 114 20878
rect 170 20822 238 20878
rect 294 20822 362 20878
rect 418 20822 486 20878
rect 542 20822 610 20878
rect 666 20822 734 20878
rect 790 20822 858 20878
rect 914 20822 982 20878
rect 1038 20822 1106 20878
rect 1162 20822 1230 20878
rect 1286 20822 1354 20878
rect 1410 20822 1478 20878
rect 1534 20822 1602 20878
rect 1658 20822 1726 20878
rect 1782 20822 1850 20878
rect 1906 20822 1916 20878
rect 104 20754 1916 20822
rect 104 20698 114 20754
rect 170 20698 238 20754
rect 294 20698 362 20754
rect 418 20698 486 20754
rect 542 20698 610 20754
rect 666 20698 734 20754
rect 790 20698 858 20754
rect 914 20698 982 20754
rect 1038 20698 1106 20754
rect 1162 20698 1230 20754
rect 1286 20698 1354 20754
rect 1410 20698 1478 20754
rect 1534 20698 1602 20754
rect 1658 20698 1726 20754
rect 1782 20698 1850 20754
rect 1906 20698 1916 20754
rect 104 20630 1916 20698
rect 104 20574 114 20630
rect 170 20574 238 20630
rect 294 20574 362 20630
rect 418 20574 486 20630
rect 542 20574 610 20630
rect 666 20574 734 20630
rect 790 20574 858 20630
rect 914 20574 982 20630
rect 1038 20574 1106 20630
rect 1162 20574 1230 20630
rect 1286 20574 1354 20630
rect 1410 20574 1478 20630
rect 1534 20574 1602 20630
rect 1658 20574 1726 20630
rect 1782 20574 1850 20630
rect 1906 20574 1916 20630
rect 104 20564 1916 20574
rect 104 20023 1916 20033
rect 104 19967 114 20023
rect 170 19967 238 20023
rect 294 19967 362 20023
rect 418 19967 486 20023
rect 542 19967 610 20023
rect 666 19967 734 20023
rect 790 19967 858 20023
rect 914 19967 982 20023
rect 1038 19967 1106 20023
rect 1162 19967 1230 20023
rect 1286 19967 1354 20023
rect 1410 19967 1478 20023
rect 1534 19967 1602 20023
rect 1658 19967 1726 20023
rect 1782 19967 1850 20023
rect 1906 19967 1916 20023
rect 104 19899 1916 19967
rect 104 19843 114 19899
rect 170 19843 238 19899
rect 294 19843 362 19899
rect 418 19843 486 19899
rect 542 19843 610 19899
rect 666 19843 734 19899
rect 790 19843 858 19899
rect 914 19843 982 19899
rect 1038 19843 1106 19899
rect 1162 19843 1230 19899
rect 1286 19843 1354 19899
rect 1410 19843 1478 19899
rect 1534 19843 1602 19899
rect 1658 19843 1726 19899
rect 1782 19843 1850 19899
rect 1906 19843 1916 19899
rect 104 19775 1916 19843
rect 104 19719 114 19775
rect 170 19719 238 19775
rect 294 19719 362 19775
rect 418 19719 486 19775
rect 542 19719 610 19775
rect 666 19719 734 19775
rect 790 19719 858 19775
rect 914 19719 982 19775
rect 1038 19719 1106 19775
rect 1162 19719 1230 19775
rect 1286 19719 1354 19775
rect 1410 19719 1478 19775
rect 1534 19719 1602 19775
rect 1658 19719 1726 19775
rect 1782 19719 1850 19775
rect 1906 19719 1916 19775
rect 104 19651 1916 19719
rect 104 19595 114 19651
rect 170 19595 238 19651
rect 294 19595 362 19651
rect 418 19595 486 19651
rect 542 19595 610 19651
rect 666 19595 734 19651
rect 790 19595 858 19651
rect 914 19595 982 19651
rect 1038 19595 1106 19651
rect 1162 19595 1230 19651
rect 1286 19595 1354 19651
rect 1410 19595 1478 19651
rect 1534 19595 1602 19651
rect 1658 19595 1726 19651
rect 1782 19595 1850 19651
rect 1906 19595 1916 19651
rect 104 19527 1916 19595
rect 104 19471 114 19527
rect 170 19471 238 19527
rect 294 19471 362 19527
rect 418 19471 486 19527
rect 542 19471 610 19527
rect 666 19471 734 19527
rect 790 19471 858 19527
rect 914 19471 982 19527
rect 1038 19471 1106 19527
rect 1162 19471 1230 19527
rect 1286 19471 1354 19527
rect 1410 19471 1478 19527
rect 1534 19471 1602 19527
rect 1658 19471 1726 19527
rect 1782 19471 1850 19527
rect 1906 19471 1916 19527
rect 104 19403 1916 19471
rect 104 19347 114 19403
rect 170 19347 238 19403
rect 294 19347 362 19403
rect 418 19347 486 19403
rect 542 19347 610 19403
rect 666 19347 734 19403
rect 790 19347 858 19403
rect 914 19347 982 19403
rect 1038 19347 1106 19403
rect 1162 19347 1230 19403
rect 1286 19347 1354 19403
rect 1410 19347 1478 19403
rect 1534 19347 1602 19403
rect 1658 19347 1726 19403
rect 1782 19347 1850 19403
rect 1906 19347 1916 19403
rect 104 19279 1916 19347
rect 104 19223 114 19279
rect 170 19223 238 19279
rect 294 19223 362 19279
rect 418 19223 486 19279
rect 542 19223 610 19279
rect 666 19223 734 19279
rect 790 19223 858 19279
rect 914 19223 982 19279
rect 1038 19223 1106 19279
rect 1162 19223 1230 19279
rect 1286 19223 1354 19279
rect 1410 19223 1478 19279
rect 1534 19223 1602 19279
rect 1658 19223 1726 19279
rect 1782 19223 1850 19279
rect 1906 19223 1916 19279
rect 104 19155 1916 19223
rect 104 19099 114 19155
rect 170 19099 238 19155
rect 294 19099 362 19155
rect 418 19099 486 19155
rect 542 19099 610 19155
rect 666 19099 734 19155
rect 790 19099 858 19155
rect 914 19099 982 19155
rect 1038 19099 1106 19155
rect 1162 19099 1230 19155
rect 1286 19099 1354 19155
rect 1410 19099 1478 19155
rect 1534 19099 1602 19155
rect 1658 19099 1726 19155
rect 1782 19099 1850 19155
rect 1906 19099 1916 19155
rect 104 19031 1916 19099
rect 104 18975 114 19031
rect 170 18975 238 19031
rect 294 18975 362 19031
rect 418 18975 486 19031
rect 542 18975 610 19031
rect 666 18975 734 19031
rect 790 18975 858 19031
rect 914 18975 982 19031
rect 1038 18975 1106 19031
rect 1162 18975 1230 19031
rect 1286 18975 1354 19031
rect 1410 18975 1478 19031
rect 1534 18975 1602 19031
rect 1658 18975 1726 19031
rect 1782 18975 1850 19031
rect 1906 18975 1916 19031
rect 104 18907 1916 18975
rect 104 18851 114 18907
rect 170 18851 238 18907
rect 294 18851 362 18907
rect 418 18851 486 18907
rect 542 18851 610 18907
rect 666 18851 734 18907
rect 790 18851 858 18907
rect 914 18851 982 18907
rect 1038 18851 1106 18907
rect 1162 18851 1230 18907
rect 1286 18851 1354 18907
rect 1410 18851 1478 18907
rect 1534 18851 1602 18907
rect 1658 18851 1726 18907
rect 1782 18851 1850 18907
rect 1906 18851 1916 18907
rect 104 18783 1916 18851
rect 104 18727 114 18783
rect 170 18727 238 18783
rect 294 18727 362 18783
rect 418 18727 486 18783
rect 542 18727 610 18783
rect 666 18727 734 18783
rect 790 18727 858 18783
rect 914 18727 982 18783
rect 1038 18727 1106 18783
rect 1162 18727 1230 18783
rect 1286 18727 1354 18783
rect 1410 18727 1478 18783
rect 1534 18727 1602 18783
rect 1658 18727 1726 18783
rect 1782 18727 1850 18783
rect 1906 18727 1916 18783
rect 104 18659 1916 18727
rect 104 18603 114 18659
rect 170 18603 238 18659
rect 294 18603 362 18659
rect 418 18603 486 18659
rect 542 18603 610 18659
rect 666 18603 734 18659
rect 790 18603 858 18659
rect 914 18603 982 18659
rect 1038 18603 1106 18659
rect 1162 18603 1230 18659
rect 1286 18603 1354 18659
rect 1410 18603 1478 18659
rect 1534 18603 1602 18659
rect 1658 18603 1726 18659
rect 1782 18603 1850 18659
rect 1906 18603 1916 18659
rect 104 18535 1916 18603
rect 104 18479 114 18535
rect 170 18479 238 18535
rect 294 18479 362 18535
rect 418 18479 486 18535
rect 542 18479 610 18535
rect 666 18479 734 18535
rect 790 18479 858 18535
rect 914 18479 982 18535
rect 1038 18479 1106 18535
rect 1162 18479 1230 18535
rect 1286 18479 1354 18535
rect 1410 18479 1478 18535
rect 1534 18479 1602 18535
rect 1658 18479 1726 18535
rect 1782 18479 1850 18535
rect 1906 18479 1916 18535
rect 104 18411 1916 18479
rect 104 18355 114 18411
rect 170 18355 238 18411
rect 294 18355 362 18411
rect 418 18355 486 18411
rect 542 18355 610 18411
rect 666 18355 734 18411
rect 790 18355 858 18411
rect 914 18355 982 18411
rect 1038 18355 1106 18411
rect 1162 18355 1230 18411
rect 1286 18355 1354 18411
rect 1410 18355 1478 18411
rect 1534 18355 1602 18411
rect 1658 18355 1726 18411
rect 1782 18355 1850 18411
rect 1906 18355 1916 18411
rect 104 18287 1916 18355
rect 104 18231 114 18287
rect 170 18231 238 18287
rect 294 18231 362 18287
rect 418 18231 486 18287
rect 542 18231 610 18287
rect 666 18231 734 18287
rect 790 18231 858 18287
rect 914 18231 982 18287
rect 1038 18231 1106 18287
rect 1162 18231 1230 18287
rect 1286 18231 1354 18287
rect 1410 18231 1478 18287
rect 1534 18231 1602 18287
rect 1658 18231 1726 18287
rect 1782 18231 1850 18287
rect 1906 18231 1916 18287
rect 104 18163 1916 18231
rect 104 18107 114 18163
rect 170 18107 238 18163
rect 294 18107 362 18163
rect 418 18107 486 18163
rect 542 18107 610 18163
rect 666 18107 734 18163
rect 790 18107 858 18163
rect 914 18107 982 18163
rect 1038 18107 1106 18163
rect 1162 18107 1230 18163
rect 1286 18107 1354 18163
rect 1410 18107 1478 18163
rect 1534 18107 1602 18163
rect 1658 18107 1726 18163
rect 1782 18107 1850 18163
rect 1906 18107 1916 18163
rect 104 18039 1916 18107
rect 104 17983 114 18039
rect 170 17983 238 18039
rect 294 17983 362 18039
rect 418 17983 486 18039
rect 542 17983 610 18039
rect 666 17983 734 18039
rect 790 17983 858 18039
rect 914 17983 982 18039
rect 1038 17983 1106 18039
rect 1162 17983 1230 18039
rect 1286 17983 1354 18039
rect 1410 17983 1478 18039
rect 1534 17983 1602 18039
rect 1658 17983 1726 18039
rect 1782 17983 1850 18039
rect 1906 17983 1916 18039
rect 104 17915 1916 17983
rect 104 17859 114 17915
rect 170 17859 238 17915
rect 294 17859 362 17915
rect 418 17859 486 17915
rect 542 17859 610 17915
rect 666 17859 734 17915
rect 790 17859 858 17915
rect 914 17859 982 17915
rect 1038 17859 1106 17915
rect 1162 17859 1230 17915
rect 1286 17859 1354 17915
rect 1410 17859 1478 17915
rect 1534 17859 1602 17915
rect 1658 17859 1726 17915
rect 1782 17859 1850 17915
rect 1906 17859 1916 17915
rect 104 17791 1916 17859
rect 104 17735 114 17791
rect 170 17735 238 17791
rect 294 17735 362 17791
rect 418 17735 486 17791
rect 542 17735 610 17791
rect 666 17735 734 17791
rect 790 17735 858 17791
rect 914 17735 982 17791
rect 1038 17735 1106 17791
rect 1162 17735 1230 17791
rect 1286 17735 1354 17791
rect 1410 17735 1478 17791
rect 1534 17735 1602 17791
rect 1658 17735 1726 17791
rect 1782 17735 1850 17791
rect 1906 17735 1916 17791
rect 104 17667 1916 17735
rect 104 17611 114 17667
rect 170 17611 238 17667
rect 294 17611 362 17667
rect 418 17611 486 17667
rect 542 17611 610 17667
rect 666 17611 734 17667
rect 790 17611 858 17667
rect 914 17611 982 17667
rect 1038 17611 1106 17667
rect 1162 17611 1230 17667
rect 1286 17611 1354 17667
rect 1410 17611 1478 17667
rect 1534 17611 1602 17667
rect 1658 17611 1726 17667
rect 1782 17611 1850 17667
rect 1906 17611 1916 17667
rect 104 17543 1916 17611
rect 104 17487 114 17543
rect 170 17487 238 17543
rect 294 17487 362 17543
rect 418 17487 486 17543
rect 542 17487 610 17543
rect 666 17487 734 17543
rect 790 17487 858 17543
rect 914 17487 982 17543
rect 1038 17487 1106 17543
rect 1162 17487 1230 17543
rect 1286 17487 1354 17543
rect 1410 17487 1478 17543
rect 1534 17487 1602 17543
rect 1658 17487 1726 17543
rect 1782 17487 1850 17543
rect 1906 17487 1916 17543
rect 104 17419 1916 17487
rect 104 17363 114 17419
rect 170 17363 238 17419
rect 294 17363 362 17419
rect 418 17363 486 17419
rect 542 17363 610 17419
rect 666 17363 734 17419
rect 790 17363 858 17419
rect 914 17363 982 17419
rect 1038 17363 1106 17419
rect 1162 17363 1230 17419
rect 1286 17363 1354 17419
rect 1410 17363 1478 17419
rect 1534 17363 1602 17419
rect 1658 17363 1726 17419
rect 1782 17363 1850 17419
rect 1906 17363 1916 17419
rect 104 17353 1916 17363
rect 104 16852 1916 16862
rect 104 16796 114 16852
rect 170 16796 238 16852
rect 294 16796 362 16852
rect 418 16796 486 16852
rect 542 16796 610 16852
rect 666 16796 734 16852
rect 790 16796 858 16852
rect 914 16796 982 16852
rect 1038 16796 1106 16852
rect 1162 16796 1230 16852
rect 1286 16796 1354 16852
rect 1410 16796 1478 16852
rect 1534 16796 1602 16852
rect 1658 16796 1726 16852
rect 1782 16796 1850 16852
rect 1906 16796 1916 16852
rect 104 16728 1916 16796
rect 104 16672 114 16728
rect 170 16672 238 16728
rect 294 16672 362 16728
rect 418 16672 486 16728
rect 542 16672 610 16728
rect 666 16672 734 16728
rect 790 16672 858 16728
rect 914 16672 982 16728
rect 1038 16672 1106 16728
rect 1162 16672 1230 16728
rect 1286 16672 1354 16728
rect 1410 16672 1478 16728
rect 1534 16672 1602 16728
rect 1658 16672 1726 16728
rect 1782 16672 1850 16728
rect 1906 16672 1916 16728
rect 104 16604 1916 16672
rect 104 16548 114 16604
rect 170 16548 238 16604
rect 294 16548 362 16604
rect 418 16548 486 16604
rect 542 16548 610 16604
rect 666 16548 734 16604
rect 790 16548 858 16604
rect 914 16548 982 16604
rect 1038 16548 1106 16604
rect 1162 16548 1230 16604
rect 1286 16548 1354 16604
rect 1410 16548 1478 16604
rect 1534 16548 1602 16604
rect 1658 16548 1726 16604
rect 1782 16548 1850 16604
rect 1906 16548 1916 16604
rect 104 16480 1916 16548
rect 104 16424 114 16480
rect 170 16424 238 16480
rect 294 16424 362 16480
rect 418 16424 486 16480
rect 542 16424 610 16480
rect 666 16424 734 16480
rect 790 16424 858 16480
rect 914 16424 982 16480
rect 1038 16424 1106 16480
rect 1162 16424 1230 16480
rect 1286 16424 1354 16480
rect 1410 16424 1478 16480
rect 1534 16424 1602 16480
rect 1658 16424 1726 16480
rect 1782 16424 1850 16480
rect 1906 16424 1916 16480
rect 104 16356 1916 16424
rect 104 16300 114 16356
rect 170 16300 238 16356
rect 294 16300 362 16356
rect 418 16300 486 16356
rect 542 16300 610 16356
rect 666 16300 734 16356
rect 790 16300 858 16356
rect 914 16300 982 16356
rect 1038 16300 1106 16356
rect 1162 16300 1230 16356
rect 1286 16300 1354 16356
rect 1410 16300 1478 16356
rect 1534 16300 1602 16356
rect 1658 16300 1726 16356
rect 1782 16300 1850 16356
rect 1906 16300 1916 16356
rect 104 16232 1916 16300
rect 104 16176 114 16232
rect 170 16176 238 16232
rect 294 16176 362 16232
rect 418 16176 486 16232
rect 542 16176 610 16232
rect 666 16176 734 16232
rect 790 16176 858 16232
rect 914 16176 982 16232
rect 1038 16176 1106 16232
rect 1162 16176 1230 16232
rect 1286 16176 1354 16232
rect 1410 16176 1478 16232
rect 1534 16176 1602 16232
rect 1658 16176 1726 16232
rect 1782 16176 1850 16232
rect 1906 16176 1916 16232
rect 104 16108 1916 16176
rect 104 16052 114 16108
rect 170 16052 238 16108
rect 294 16052 362 16108
rect 418 16052 486 16108
rect 542 16052 610 16108
rect 666 16052 734 16108
rect 790 16052 858 16108
rect 914 16052 982 16108
rect 1038 16052 1106 16108
rect 1162 16052 1230 16108
rect 1286 16052 1354 16108
rect 1410 16052 1478 16108
rect 1534 16052 1602 16108
rect 1658 16052 1726 16108
rect 1782 16052 1850 16108
rect 1906 16052 1916 16108
rect 104 15984 1916 16052
rect 104 15928 114 15984
rect 170 15928 238 15984
rect 294 15928 362 15984
rect 418 15928 486 15984
rect 542 15928 610 15984
rect 666 15928 734 15984
rect 790 15928 858 15984
rect 914 15928 982 15984
rect 1038 15928 1106 15984
rect 1162 15928 1230 15984
rect 1286 15928 1354 15984
rect 1410 15928 1478 15984
rect 1534 15928 1602 15984
rect 1658 15928 1726 15984
rect 1782 15928 1850 15984
rect 1906 15928 1916 15984
rect 104 15860 1916 15928
rect 104 15804 114 15860
rect 170 15804 238 15860
rect 294 15804 362 15860
rect 418 15804 486 15860
rect 542 15804 610 15860
rect 666 15804 734 15860
rect 790 15804 858 15860
rect 914 15804 982 15860
rect 1038 15804 1106 15860
rect 1162 15804 1230 15860
rect 1286 15804 1354 15860
rect 1410 15804 1478 15860
rect 1534 15804 1602 15860
rect 1658 15804 1726 15860
rect 1782 15804 1850 15860
rect 1906 15804 1916 15860
rect 104 15736 1916 15804
rect 104 15680 114 15736
rect 170 15680 238 15736
rect 294 15680 362 15736
rect 418 15680 486 15736
rect 542 15680 610 15736
rect 666 15680 734 15736
rect 790 15680 858 15736
rect 914 15680 982 15736
rect 1038 15680 1106 15736
rect 1162 15680 1230 15736
rect 1286 15680 1354 15736
rect 1410 15680 1478 15736
rect 1534 15680 1602 15736
rect 1658 15680 1726 15736
rect 1782 15680 1850 15736
rect 1906 15680 1916 15736
rect 104 15612 1916 15680
rect 104 15556 114 15612
rect 170 15556 238 15612
rect 294 15556 362 15612
rect 418 15556 486 15612
rect 542 15556 610 15612
rect 666 15556 734 15612
rect 790 15556 858 15612
rect 914 15556 982 15612
rect 1038 15556 1106 15612
rect 1162 15556 1230 15612
rect 1286 15556 1354 15612
rect 1410 15556 1478 15612
rect 1534 15556 1602 15612
rect 1658 15556 1726 15612
rect 1782 15556 1850 15612
rect 1906 15556 1916 15612
rect 104 15488 1916 15556
rect 104 15432 114 15488
rect 170 15432 238 15488
rect 294 15432 362 15488
rect 418 15432 486 15488
rect 542 15432 610 15488
rect 666 15432 734 15488
rect 790 15432 858 15488
rect 914 15432 982 15488
rect 1038 15432 1106 15488
rect 1162 15432 1230 15488
rect 1286 15432 1354 15488
rect 1410 15432 1478 15488
rect 1534 15432 1602 15488
rect 1658 15432 1726 15488
rect 1782 15432 1850 15488
rect 1906 15432 1916 15488
rect 104 15364 1916 15432
rect 104 15308 114 15364
rect 170 15308 238 15364
rect 294 15308 362 15364
rect 418 15308 486 15364
rect 542 15308 610 15364
rect 666 15308 734 15364
rect 790 15308 858 15364
rect 914 15308 982 15364
rect 1038 15308 1106 15364
rect 1162 15308 1230 15364
rect 1286 15308 1354 15364
rect 1410 15308 1478 15364
rect 1534 15308 1602 15364
rect 1658 15308 1726 15364
rect 1782 15308 1850 15364
rect 1906 15308 1916 15364
rect 104 15240 1916 15308
rect 104 15184 114 15240
rect 170 15184 238 15240
rect 294 15184 362 15240
rect 418 15184 486 15240
rect 542 15184 610 15240
rect 666 15184 734 15240
rect 790 15184 858 15240
rect 914 15184 982 15240
rect 1038 15184 1106 15240
rect 1162 15184 1230 15240
rect 1286 15184 1354 15240
rect 1410 15184 1478 15240
rect 1534 15184 1602 15240
rect 1658 15184 1726 15240
rect 1782 15184 1850 15240
rect 1906 15184 1916 15240
rect 104 15116 1916 15184
rect 104 15060 114 15116
rect 170 15060 238 15116
rect 294 15060 362 15116
rect 418 15060 486 15116
rect 542 15060 610 15116
rect 666 15060 734 15116
rect 790 15060 858 15116
rect 914 15060 982 15116
rect 1038 15060 1106 15116
rect 1162 15060 1230 15116
rect 1286 15060 1354 15116
rect 1410 15060 1478 15116
rect 1534 15060 1602 15116
rect 1658 15060 1726 15116
rect 1782 15060 1850 15116
rect 1906 15060 1916 15116
rect 104 14992 1916 15060
rect 104 14936 114 14992
rect 170 14936 238 14992
rect 294 14936 362 14992
rect 418 14936 486 14992
rect 542 14936 610 14992
rect 666 14936 734 14992
rect 790 14936 858 14992
rect 914 14936 982 14992
rect 1038 14936 1106 14992
rect 1162 14936 1230 14992
rect 1286 14936 1354 14992
rect 1410 14936 1478 14992
rect 1534 14936 1602 14992
rect 1658 14936 1726 14992
rect 1782 14936 1850 14992
rect 1906 14936 1916 14992
rect 104 14868 1916 14936
rect 104 14812 114 14868
rect 170 14812 238 14868
rect 294 14812 362 14868
rect 418 14812 486 14868
rect 542 14812 610 14868
rect 666 14812 734 14868
rect 790 14812 858 14868
rect 914 14812 982 14868
rect 1038 14812 1106 14868
rect 1162 14812 1230 14868
rect 1286 14812 1354 14868
rect 1410 14812 1478 14868
rect 1534 14812 1602 14868
rect 1658 14812 1726 14868
rect 1782 14812 1850 14868
rect 1906 14812 1916 14868
rect 104 14744 1916 14812
rect 104 14688 114 14744
rect 170 14688 238 14744
rect 294 14688 362 14744
rect 418 14688 486 14744
rect 542 14688 610 14744
rect 666 14688 734 14744
rect 790 14688 858 14744
rect 914 14688 982 14744
rect 1038 14688 1106 14744
rect 1162 14688 1230 14744
rect 1286 14688 1354 14744
rect 1410 14688 1478 14744
rect 1534 14688 1602 14744
rect 1658 14688 1726 14744
rect 1782 14688 1850 14744
rect 1906 14688 1916 14744
rect 104 14620 1916 14688
rect 104 14564 114 14620
rect 170 14564 238 14620
rect 294 14564 362 14620
rect 418 14564 486 14620
rect 542 14564 610 14620
rect 666 14564 734 14620
rect 790 14564 858 14620
rect 914 14564 982 14620
rect 1038 14564 1106 14620
rect 1162 14564 1230 14620
rect 1286 14564 1354 14620
rect 1410 14564 1478 14620
rect 1534 14564 1602 14620
rect 1658 14564 1726 14620
rect 1782 14564 1850 14620
rect 1906 14564 1916 14620
rect 104 14496 1916 14564
rect 104 14440 114 14496
rect 170 14440 238 14496
rect 294 14440 362 14496
rect 418 14440 486 14496
rect 542 14440 610 14496
rect 666 14440 734 14496
rect 790 14440 858 14496
rect 914 14440 982 14496
rect 1038 14440 1106 14496
rect 1162 14440 1230 14496
rect 1286 14440 1354 14496
rect 1410 14440 1478 14496
rect 1534 14440 1602 14496
rect 1658 14440 1726 14496
rect 1782 14440 1850 14496
rect 1906 14440 1916 14496
rect 104 14372 1916 14440
rect 104 14316 114 14372
rect 170 14316 238 14372
rect 294 14316 362 14372
rect 418 14316 486 14372
rect 542 14316 610 14372
rect 666 14316 734 14372
rect 790 14316 858 14372
rect 914 14316 982 14372
rect 1038 14316 1106 14372
rect 1162 14316 1230 14372
rect 1286 14316 1354 14372
rect 1410 14316 1478 14372
rect 1534 14316 1602 14372
rect 1658 14316 1726 14372
rect 1782 14316 1850 14372
rect 1906 14316 1916 14372
rect 104 14248 1916 14316
rect 104 14192 114 14248
rect 170 14192 238 14248
rect 294 14192 362 14248
rect 418 14192 486 14248
rect 542 14192 610 14248
rect 666 14192 734 14248
rect 790 14192 858 14248
rect 914 14192 982 14248
rect 1038 14192 1106 14248
rect 1162 14192 1230 14248
rect 1286 14192 1354 14248
rect 1410 14192 1478 14248
rect 1534 14192 1602 14248
rect 1658 14192 1726 14248
rect 1782 14192 1850 14248
rect 1906 14192 1916 14248
rect 104 14182 1916 14192
<< via3 >>
rect 114 69568 170 69624
rect 238 69568 294 69624
rect 362 69568 418 69624
rect 486 69568 542 69624
rect 610 69568 666 69624
rect 734 69568 790 69624
rect 858 69568 914 69624
rect 982 69568 1038 69624
rect 1106 69568 1162 69624
rect 1230 69568 1286 69624
rect 1354 69568 1410 69624
rect 1478 69568 1534 69624
rect 1602 69568 1658 69624
rect 1726 69568 1782 69624
rect 1850 69568 1906 69624
rect 114 69444 170 69500
rect 238 69444 294 69500
rect 362 69444 418 69500
rect 486 69444 542 69500
rect 610 69444 666 69500
rect 734 69444 790 69500
rect 858 69444 914 69500
rect 982 69444 1038 69500
rect 1106 69444 1162 69500
rect 1230 69444 1286 69500
rect 1354 69444 1410 69500
rect 1478 69444 1534 69500
rect 1602 69444 1658 69500
rect 1726 69444 1782 69500
rect 1850 69444 1906 69500
rect 114 69320 170 69376
rect 238 69320 294 69376
rect 362 69320 418 69376
rect 486 69320 542 69376
rect 610 69320 666 69376
rect 734 69320 790 69376
rect 858 69320 914 69376
rect 982 69320 1038 69376
rect 1106 69320 1162 69376
rect 1230 69320 1286 69376
rect 1354 69320 1410 69376
rect 1478 69320 1534 69376
rect 1602 69320 1658 69376
rect 1726 69320 1782 69376
rect 1850 69320 1906 69376
rect 114 69196 170 69252
rect 238 69196 294 69252
rect 362 69196 418 69252
rect 486 69196 542 69252
rect 610 69196 666 69252
rect 734 69196 790 69252
rect 858 69196 914 69252
rect 982 69196 1038 69252
rect 1106 69196 1162 69252
rect 1230 69196 1286 69252
rect 1354 69196 1410 69252
rect 1478 69196 1534 69252
rect 1602 69196 1658 69252
rect 1726 69196 1782 69252
rect 1850 69196 1906 69252
rect 114 69072 170 69128
rect 238 69072 294 69128
rect 362 69072 418 69128
rect 486 69072 542 69128
rect 610 69072 666 69128
rect 734 69072 790 69128
rect 858 69072 914 69128
rect 982 69072 1038 69128
rect 1106 69072 1162 69128
rect 1230 69072 1286 69128
rect 1354 69072 1410 69128
rect 1478 69072 1534 69128
rect 1602 69072 1658 69128
rect 1726 69072 1782 69128
rect 1850 69072 1906 69128
rect 114 68948 170 69004
rect 238 68948 294 69004
rect 362 68948 418 69004
rect 486 68948 542 69004
rect 610 68948 666 69004
rect 734 68948 790 69004
rect 858 68948 914 69004
rect 982 68948 1038 69004
rect 1106 68948 1162 69004
rect 1230 68948 1286 69004
rect 1354 68948 1410 69004
rect 1478 68948 1534 69004
rect 1602 68948 1658 69004
rect 1726 68948 1782 69004
rect 1850 68948 1906 69004
rect 114 68824 170 68880
rect 238 68824 294 68880
rect 362 68824 418 68880
rect 486 68824 542 68880
rect 610 68824 666 68880
rect 734 68824 790 68880
rect 858 68824 914 68880
rect 982 68824 1038 68880
rect 1106 68824 1162 68880
rect 1230 68824 1286 68880
rect 1354 68824 1410 68880
rect 1478 68824 1534 68880
rect 1602 68824 1658 68880
rect 1726 68824 1782 68880
rect 1850 68824 1906 68880
rect 114 68700 170 68756
rect 238 68700 294 68756
rect 362 68700 418 68756
rect 486 68700 542 68756
rect 610 68700 666 68756
rect 734 68700 790 68756
rect 858 68700 914 68756
rect 982 68700 1038 68756
rect 1106 68700 1162 68756
rect 1230 68700 1286 68756
rect 1354 68700 1410 68756
rect 1478 68700 1534 68756
rect 1602 68700 1658 68756
rect 1726 68700 1782 68756
rect 1850 68700 1906 68756
rect 114 68576 170 68632
rect 238 68576 294 68632
rect 362 68576 418 68632
rect 486 68576 542 68632
rect 610 68576 666 68632
rect 734 68576 790 68632
rect 858 68576 914 68632
rect 982 68576 1038 68632
rect 1106 68576 1162 68632
rect 1230 68576 1286 68632
rect 1354 68576 1410 68632
rect 1478 68576 1534 68632
rect 1602 68576 1658 68632
rect 1726 68576 1782 68632
rect 1850 68576 1906 68632
rect 114 68452 170 68508
rect 238 68452 294 68508
rect 362 68452 418 68508
rect 486 68452 542 68508
rect 610 68452 666 68508
rect 734 68452 790 68508
rect 858 68452 914 68508
rect 982 68452 1038 68508
rect 1106 68452 1162 68508
rect 1230 68452 1286 68508
rect 1354 68452 1410 68508
rect 1478 68452 1534 68508
rect 1602 68452 1658 68508
rect 1726 68452 1782 68508
rect 1850 68452 1906 68508
rect 114 68038 170 68094
rect 238 68038 294 68094
rect 362 68038 418 68094
rect 486 68038 542 68094
rect 610 68038 666 68094
rect 734 68038 790 68094
rect 858 68038 914 68094
rect 982 68038 1038 68094
rect 1106 68038 1162 68094
rect 1230 68038 1286 68094
rect 1354 68038 1410 68094
rect 1478 68038 1534 68094
rect 1602 68038 1658 68094
rect 1726 68038 1782 68094
rect 1850 68038 1906 68094
rect 114 67914 170 67970
rect 238 67914 294 67970
rect 362 67914 418 67970
rect 486 67914 542 67970
rect 610 67914 666 67970
rect 734 67914 790 67970
rect 858 67914 914 67970
rect 982 67914 1038 67970
rect 1106 67914 1162 67970
rect 1230 67914 1286 67970
rect 1354 67914 1410 67970
rect 1478 67914 1534 67970
rect 1602 67914 1658 67970
rect 1726 67914 1782 67970
rect 1850 67914 1906 67970
rect 114 67790 170 67846
rect 238 67790 294 67846
rect 362 67790 418 67846
rect 486 67790 542 67846
rect 610 67790 666 67846
rect 734 67790 790 67846
rect 858 67790 914 67846
rect 982 67790 1038 67846
rect 1106 67790 1162 67846
rect 1230 67790 1286 67846
rect 1354 67790 1410 67846
rect 1478 67790 1534 67846
rect 1602 67790 1658 67846
rect 1726 67790 1782 67846
rect 1850 67790 1906 67846
rect 114 67666 170 67722
rect 238 67666 294 67722
rect 362 67666 418 67722
rect 486 67666 542 67722
rect 610 67666 666 67722
rect 734 67666 790 67722
rect 858 67666 914 67722
rect 982 67666 1038 67722
rect 1106 67666 1162 67722
rect 1230 67666 1286 67722
rect 1354 67666 1410 67722
rect 1478 67666 1534 67722
rect 1602 67666 1658 67722
rect 1726 67666 1782 67722
rect 1850 67666 1906 67722
rect 114 67542 170 67598
rect 238 67542 294 67598
rect 362 67542 418 67598
rect 486 67542 542 67598
rect 610 67542 666 67598
rect 734 67542 790 67598
rect 858 67542 914 67598
rect 982 67542 1038 67598
rect 1106 67542 1162 67598
rect 1230 67542 1286 67598
rect 1354 67542 1410 67598
rect 1478 67542 1534 67598
rect 1602 67542 1658 67598
rect 1726 67542 1782 67598
rect 1850 67542 1906 67598
rect 114 67418 170 67474
rect 238 67418 294 67474
rect 362 67418 418 67474
rect 486 67418 542 67474
rect 610 67418 666 67474
rect 734 67418 790 67474
rect 858 67418 914 67474
rect 982 67418 1038 67474
rect 1106 67418 1162 67474
rect 1230 67418 1286 67474
rect 1354 67418 1410 67474
rect 1478 67418 1534 67474
rect 1602 67418 1658 67474
rect 1726 67418 1782 67474
rect 1850 67418 1906 67474
rect 114 67294 170 67350
rect 238 67294 294 67350
rect 362 67294 418 67350
rect 486 67294 542 67350
rect 610 67294 666 67350
rect 734 67294 790 67350
rect 858 67294 914 67350
rect 982 67294 1038 67350
rect 1106 67294 1162 67350
rect 1230 67294 1286 67350
rect 1354 67294 1410 67350
rect 1478 67294 1534 67350
rect 1602 67294 1658 67350
rect 1726 67294 1782 67350
rect 1850 67294 1906 67350
rect 114 67170 170 67226
rect 238 67170 294 67226
rect 362 67170 418 67226
rect 486 67170 542 67226
rect 610 67170 666 67226
rect 734 67170 790 67226
rect 858 67170 914 67226
rect 982 67170 1038 67226
rect 1106 67170 1162 67226
rect 1230 67170 1286 67226
rect 1354 67170 1410 67226
rect 1478 67170 1534 67226
rect 1602 67170 1658 67226
rect 1726 67170 1782 67226
rect 1850 67170 1906 67226
rect 114 67046 170 67102
rect 238 67046 294 67102
rect 362 67046 418 67102
rect 486 67046 542 67102
rect 610 67046 666 67102
rect 734 67046 790 67102
rect 858 67046 914 67102
rect 982 67046 1038 67102
rect 1106 67046 1162 67102
rect 1230 67046 1286 67102
rect 1354 67046 1410 67102
rect 1478 67046 1534 67102
rect 1602 67046 1658 67102
rect 1726 67046 1782 67102
rect 1850 67046 1906 67102
rect 114 66922 170 66978
rect 238 66922 294 66978
rect 362 66922 418 66978
rect 486 66922 542 66978
rect 610 66922 666 66978
rect 734 66922 790 66978
rect 858 66922 914 66978
rect 982 66922 1038 66978
rect 1106 66922 1162 66978
rect 1230 66922 1286 66978
rect 1354 66922 1410 66978
rect 1478 66922 1534 66978
rect 1602 66922 1658 66978
rect 1726 66922 1782 66978
rect 1850 66922 1906 66978
rect 114 66428 170 66484
rect 238 66428 294 66484
rect 362 66428 418 66484
rect 486 66428 542 66484
rect 610 66428 666 66484
rect 734 66428 790 66484
rect 858 66428 914 66484
rect 982 66428 1038 66484
rect 1106 66428 1162 66484
rect 1230 66428 1286 66484
rect 1354 66428 1410 66484
rect 1478 66428 1534 66484
rect 1602 66428 1658 66484
rect 1726 66428 1782 66484
rect 1850 66428 1906 66484
rect 114 66304 170 66360
rect 238 66304 294 66360
rect 362 66304 418 66360
rect 486 66304 542 66360
rect 610 66304 666 66360
rect 734 66304 790 66360
rect 858 66304 914 66360
rect 982 66304 1038 66360
rect 1106 66304 1162 66360
rect 1230 66304 1286 66360
rect 1354 66304 1410 66360
rect 1478 66304 1534 66360
rect 1602 66304 1658 66360
rect 1726 66304 1782 66360
rect 1850 66304 1906 66360
rect 114 66180 170 66236
rect 238 66180 294 66236
rect 362 66180 418 66236
rect 486 66180 542 66236
rect 610 66180 666 66236
rect 734 66180 790 66236
rect 858 66180 914 66236
rect 982 66180 1038 66236
rect 1106 66180 1162 66236
rect 1230 66180 1286 66236
rect 1354 66180 1410 66236
rect 1478 66180 1534 66236
rect 1602 66180 1658 66236
rect 1726 66180 1782 66236
rect 1850 66180 1906 66236
rect 114 66056 170 66112
rect 238 66056 294 66112
rect 362 66056 418 66112
rect 486 66056 542 66112
rect 610 66056 666 66112
rect 734 66056 790 66112
rect 858 66056 914 66112
rect 982 66056 1038 66112
rect 1106 66056 1162 66112
rect 1230 66056 1286 66112
rect 1354 66056 1410 66112
rect 1478 66056 1534 66112
rect 1602 66056 1658 66112
rect 1726 66056 1782 66112
rect 1850 66056 1906 66112
rect 114 65932 170 65988
rect 238 65932 294 65988
rect 362 65932 418 65988
rect 486 65932 542 65988
rect 610 65932 666 65988
rect 734 65932 790 65988
rect 858 65932 914 65988
rect 982 65932 1038 65988
rect 1106 65932 1162 65988
rect 1230 65932 1286 65988
rect 1354 65932 1410 65988
rect 1478 65932 1534 65988
rect 1602 65932 1658 65988
rect 1726 65932 1782 65988
rect 1850 65932 1906 65988
rect 114 65808 170 65864
rect 238 65808 294 65864
rect 362 65808 418 65864
rect 486 65808 542 65864
rect 610 65808 666 65864
rect 734 65808 790 65864
rect 858 65808 914 65864
rect 982 65808 1038 65864
rect 1106 65808 1162 65864
rect 1230 65808 1286 65864
rect 1354 65808 1410 65864
rect 1478 65808 1534 65864
rect 1602 65808 1658 65864
rect 1726 65808 1782 65864
rect 1850 65808 1906 65864
rect 114 65684 170 65740
rect 238 65684 294 65740
rect 362 65684 418 65740
rect 486 65684 542 65740
rect 610 65684 666 65740
rect 734 65684 790 65740
rect 858 65684 914 65740
rect 982 65684 1038 65740
rect 1106 65684 1162 65740
rect 1230 65684 1286 65740
rect 1354 65684 1410 65740
rect 1478 65684 1534 65740
rect 1602 65684 1658 65740
rect 1726 65684 1782 65740
rect 1850 65684 1906 65740
rect 114 65560 170 65616
rect 238 65560 294 65616
rect 362 65560 418 65616
rect 486 65560 542 65616
rect 610 65560 666 65616
rect 734 65560 790 65616
rect 858 65560 914 65616
rect 982 65560 1038 65616
rect 1106 65560 1162 65616
rect 1230 65560 1286 65616
rect 1354 65560 1410 65616
rect 1478 65560 1534 65616
rect 1602 65560 1658 65616
rect 1726 65560 1782 65616
rect 1850 65560 1906 65616
rect 114 65436 170 65492
rect 238 65436 294 65492
rect 362 65436 418 65492
rect 486 65436 542 65492
rect 610 65436 666 65492
rect 734 65436 790 65492
rect 858 65436 914 65492
rect 982 65436 1038 65492
rect 1106 65436 1162 65492
rect 1230 65436 1286 65492
rect 1354 65436 1410 65492
rect 1478 65436 1534 65492
rect 1602 65436 1658 65492
rect 1726 65436 1782 65492
rect 1850 65436 1906 65492
rect 114 65312 170 65368
rect 238 65312 294 65368
rect 362 65312 418 65368
rect 486 65312 542 65368
rect 610 65312 666 65368
rect 734 65312 790 65368
rect 858 65312 914 65368
rect 982 65312 1038 65368
rect 1106 65312 1162 65368
rect 1230 65312 1286 65368
rect 1354 65312 1410 65368
rect 1478 65312 1534 65368
rect 1602 65312 1658 65368
rect 1726 65312 1782 65368
rect 1850 65312 1906 65368
rect 114 64830 170 64886
rect 238 64830 294 64886
rect 362 64830 418 64886
rect 486 64830 542 64886
rect 610 64830 666 64886
rect 734 64830 790 64886
rect 858 64830 914 64886
rect 982 64830 1038 64886
rect 1106 64830 1162 64886
rect 1230 64830 1286 64886
rect 1354 64830 1410 64886
rect 1478 64830 1534 64886
rect 1602 64830 1658 64886
rect 1726 64830 1782 64886
rect 1850 64830 1906 64886
rect 114 64706 170 64762
rect 238 64706 294 64762
rect 362 64706 418 64762
rect 486 64706 542 64762
rect 610 64706 666 64762
rect 734 64706 790 64762
rect 858 64706 914 64762
rect 982 64706 1038 64762
rect 1106 64706 1162 64762
rect 1230 64706 1286 64762
rect 1354 64706 1410 64762
rect 1478 64706 1534 64762
rect 1602 64706 1658 64762
rect 1726 64706 1782 64762
rect 1850 64706 1906 64762
rect 114 64582 170 64638
rect 238 64582 294 64638
rect 362 64582 418 64638
rect 486 64582 542 64638
rect 610 64582 666 64638
rect 734 64582 790 64638
rect 858 64582 914 64638
rect 982 64582 1038 64638
rect 1106 64582 1162 64638
rect 1230 64582 1286 64638
rect 1354 64582 1410 64638
rect 1478 64582 1534 64638
rect 1602 64582 1658 64638
rect 1726 64582 1782 64638
rect 1850 64582 1906 64638
rect 114 64458 170 64514
rect 238 64458 294 64514
rect 362 64458 418 64514
rect 486 64458 542 64514
rect 610 64458 666 64514
rect 734 64458 790 64514
rect 858 64458 914 64514
rect 982 64458 1038 64514
rect 1106 64458 1162 64514
rect 1230 64458 1286 64514
rect 1354 64458 1410 64514
rect 1478 64458 1534 64514
rect 1602 64458 1658 64514
rect 1726 64458 1782 64514
rect 1850 64458 1906 64514
rect 114 64334 170 64390
rect 238 64334 294 64390
rect 362 64334 418 64390
rect 486 64334 542 64390
rect 610 64334 666 64390
rect 734 64334 790 64390
rect 858 64334 914 64390
rect 982 64334 1038 64390
rect 1106 64334 1162 64390
rect 1230 64334 1286 64390
rect 1354 64334 1410 64390
rect 1478 64334 1534 64390
rect 1602 64334 1658 64390
rect 1726 64334 1782 64390
rect 1850 64334 1906 64390
rect 114 64210 170 64266
rect 238 64210 294 64266
rect 362 64210 418 64266
rect 486 64210 542 64266
rect 610 64210 666 64266
rect 734 64210 790 64266
rect 858 64210 914 64266
rect 982 64210 1038 64266
rect 1106 64210 1162 64266
rect 1230 64210 1286 64266
rect 1354 64210 1410 64266
rect 1478 64210 1534 64266
rect 1602 64210 1658 64266
rect 1726 64210 1782 64266
rect 1850 64210 1906 64266
rect 114 64086 170 64142
rect 238 64086 294 64142
rect 362 64086 418 64142
rect 486 64086 542 64142
rect 610 64086 666 64142
rect 734 64086 790 64142
rect 858 64086 914 64142
rect 982 64086 1038 64142
rect 1106 64086 1162 64142
rect 1230 64086 1286 64142
rect 1354 64086 1410 64142
rect 1478 64086 1534 64142
rect 1602 64086 1658 64142
rect 1726 64086 1782 64142
rect 1850 64086 1906 64142
rect 114 63962 170 64018
rect 238 63962 294 64018
rect 362 63962 418 64018
rect 486 63962 542 64018
rect 610 63962 666 64018
rect 734 63962 790 64018
rect 858 63962 914 64018
rect 982 63962 1038 64018
rect 1106 63962 1162 64018
rect 1230 63962 1286 64018
rect 1354 63962 1410 64018
rect 1478 63962 1534 64018
rect 1602 63962 1658 64018
rect 1726 63962 1782 64018
rect 1850 63962 1906 64018
rect 114 63838 170 63894
rect 238 63838 294 63894
rect 362 63838 418 63894
rect 486 63838 542 63894
rect 610 63838 666 63894
rect 734 63838 790 63894
rect 858 63838 914 63894
rect 982 63838 1038 63894
rect 1106 63838 1162 63894
rect 1230 63838 1286 63894
rect 1354 63838 1410 63894
rect 1478 63838 1534 63894
rect 1602 63838 1658 63894
rect 1726 63838 1782 63894
rect 1850 63838 1906 63894
rect 114 63714 170 63770
rect 238 63714 294 63770
rect 362 63714 418 63770
rect 486 63714 542 63770
rect 610 63714 666 63770
rect 734 63714 790 63770
rect 858 63714 914 63770
rect 982 63714 1038 63770
rect 1106 63714 1162 63770
rect 1230 63714 1286 63770
rect 1354 63714 1410 63770
rect 1478 63714 1534 63770
rect 1602 63714 1658 63770
rect 1726 63714 1782 63770
rect 1850 63714 1906 63770
rect 114 63239 170 63295
rect 238 63239 294 63295
rect 362 63239 418 63295
rect 486 63239 542 63295
rect 610 63239 666 63295
rect 734 63239 790 63295
rect 858 63239 914 63295
rect 982 63239 1038 63295
rect 1106 63239 1162 63295
rect 1230 63239 1286 63295
rect 1354 63239 1410 63295
rect 1478 63239 1534 63295
rect 1602 63239 1658 63295
rect 1726 63239 1782 63295
rect 1850 63239 1906 63295
rect 114 63115 170 63171
rect 238 63115 294 63171
rect 362 63115 418 63171
rect 486 63115 542 63171
rect 610 63115 666 63171
rect 734 63115 790 63171
rect 858 63115 914 63171
rect 982 63115 1038 63171
rect 1106 63115 1162 63171
rect 1230 63115 1286 63171
rect 1354 63115 1410 63171
rect 1478 63115 1534 63171
rect 1602 63115 1658 63171
rect 1726 63115 1782 63171
rect 1850 63115 1906 63171
rect 114 62991 170 63047
rect 238 62991 294 63047
rect 362 62991 418 63047
rect 486 62991 542 63047
rect 610 62991 666 63047
rect 734 62991 790 63047
rect 858 62991 914 63047
rect 982 62991 1038 63047
rect 1106 62991 1162 63047
rect 1230 62991 1286 63047
rect 1354 62991 1410 63047
rect 1478 62991 1534 63047
rect 1602 62991 1658 63047
rect 1726 62991 1782 63047
rect 1850 62991 1906 63047
rect 114 62867 170 62923
rect 238 62867 294 62923
rect 362 62867 418 62923
rect 486 62867 542 62923
rect 610 62867 666 62923
rect 734 62867 790 62923
rect 858 62867 914 62923
rect 982 62867 1038 62923
rect 1106 62867 1162 62923
rect 1230 62867 1286 62923
rect 1354 62867 1410 62923
rect 1478 62867 1534 62923
rect 1602 62867 1658 62923
rect 1726 62867 1782 62923
rect 1850 62867 1906 62923
rect 114 62743 170 62799
rect 238 62743 294 62799
rect 362 62743 418 62799
rect 486 62743 542 62799
rect 610 62743 666 62799
rect 734 62743 790 62799
rect 858 62743 914 62799
rect 982 62743 1038 62799
rect 1106 62743 1162 62799
rect 1230 62743 1286 62799
rect 1354 62743 1410 62799
rect 1478 62743 1534 62799
rect 1602 62743 1658 62799
rect 1726 62743 1782 62799
rect 1850 62743 1906 62799
rect 114 62619 170 62675
rect 238 62619 294 62675
rect 362 62619 418 62675
rect 486 62619 542 62675
rect 610 62619 666 62675
rect 734 62619 790 62675
rect 858 62619 914 62675
rect 982 62619 1038 62675
rect 1106 62619 1162 62675
rect 1230 62619 1286 62675
rect 1354 62619 1410 62675
rect 1478 62619 1534 62675
rect 1602 62619 1658 62675
rect 1726 62619 1782 62675
rect 1850 62619 1906 62675
rect 114 62495 170 62551
rect 238 62495 294 62551
rect 362 62495 418 62551
rect 486 62495 542 62551
rect 610 62495 666 62551
rect 734 62495 790 62551
rect 858 62495 914 62551
rect 982 62495 1038 62551
rect 1106 62495 1162 62551
rect 1230 62495 1286 62551
rect 1354 62495 1410 62551
rect 1478 62495 1534 62551
rect 1602 62495 1658 62551
rect 1726 62495 1782 62551
rect 1850 62495 1906 62551
rect 114 62371 170 62427
rect 238 62371 294 62427
rect 362 62371 418 62427
rect 486 62371 542 62427
rect 610 62371 666 62427
rect 734 62371 790 62427
rect 858 62371 914 62427
rect 982 62371 1038 62427
rect 1106 62371 1162 62427
rect 1230 62371 1286 62427
rect 1354 62371 1410 62427
rect 1478 62371 1534 62427
rect 1602 62371 1658 62427
rect 1726 62371 1782 62427
rect 1850 62371 1906 62427
rect 114 62247 170 62303
rect 238 62247 294 62303
rect 362 62247 418 62303
rect 486 62247 542 62303
rect 610 62247 666 62303
rect 734 62247 790 62303
rect 858 62247 914 62303
rect 982 62247 1038 62303
rect 1106 62247 1162 62303
rect 1230 62247 1286 62303
rect 1354 62247 1410 62303
rect 1478 62247 1534 62303
rect 1602 62247 1658 62303
rect 1726 62247 1782 62303
rect 1850 62247 1906 62303
rect 114 62123 170 62179
rect 238 62123 294 62179
rect 362 62123 418 62179
rect 486 62123 542 62179
rect 610 62123 666 62179
rect 734 62123 790 62179
rect 858 62123 914 62179
rect 982 62123 1038 62179
rect 1106 62123 1162 62179
rect 1230 62123 1286 62179
rect 1354 62123 1410 62179
rect 1478 62123 1534 62179
rect 1602 62123 1658 62179
rect 1726 62123 1782 62179
rect 1850 62123 1906 62179
rect 114 61639 170 61695
rect 238 61639 294 61695
rect 362 61639 418 61695
rect 486 61639 542 61695
rect 610 61639 666 61695
rect 734 61639 790 61695
rect 858 61639 914 61695
rect 982 61639 1038 61695
rect 1106 61639 1162 61695
rect 1230 61639 1286 61695
rect 1354 61639 1410 61695
rect 1478 61639 1534 61695
rect 1602 61639 1658 61695
rect 1726 61639 1782 61695
rect 1850 61639 1906 61695
rect 114 61515 170 61571
rect 238 61515 294 61571
rect 362 61515 418 61571
rect 486 61515 542 61571
rect 610 61515 666 61571
rect 734 61515 790 61571
rect 858 61515 914 61571
rect 982 61515 1038 61571
rect 1106 61515 1162 61571
rect 1230 61515 1286 61571
rect 1354 61515 1410 61571
rect 1478 61515 1534 61571
rect 1602 61515 1658 61571
rect 1726 61515 1782 61571
rect 1850 61515 1906 61571
rect 114 61391 170 61447
rect 238 61391 294 61447
rect 362 61391 418 61447
rect 486 61391 542 61447
rect 610 61391 666 61447
rect 734 61391 790 61447
rect 858 61391 914 61447
rect 982 61391 1038 61447
rect 1106 61391 1162 61447
rect 1230 61391 1286 61447
rect 1354 61391 1410 61447
rect 1478 61391 1534 61447
rect 1602 61391 1658 61447
rect 1726 61391 1782 61447
rect 1850 61391 1906 61447
rect 114 61267 170 61323
rect 238 61267 294 61323
rect 362 61267 418 61323
rect 486 61267 542 61323
rect 610 61267 666 61323
rect 734 61267 790 61323
rect 858 61267 914 61323
rect 982 61267 1038 61323
rect 1106 61267 1162 61323
rect 1230 61267 1286 61323
rect 1354 61267 1410 61323
rect 1478 61267 1534 61323
rect 1602 61267 1658 61323
rect 1726 61267 1782 61323
rect 1850 61267 1906 61323
rect 114 61143 170 61199
rect 238 61143 294 61199
rect 362 61143 418 61199
rect 486 61143 542 61199
rect 610 61143 666 61199
rect 734 61143 790 61199
rect 858 61143 914 61199
rect 982 61143 1038 61199
rect 1106 61143 1162 61199
rect 1230 61143 1286 61199
rect 1354 61143 1410 61199
rect 1478 61143 1534 61199
rect 1602 61143 1658 61199
rect 1726 61143 1782 61199
rect 1850 61143 1906 61199
rect 114 61019 170 61075
rect 238 61019 294 61075
rect 362 61019 418 61075
rect 486 61019 542 61075
rect 610 61019 666 61075
rect 734 61019 790 61075
rect 858 61019 914 61075
rect 982 61019 1038 61075
rect 1106 61019 1162 61075
rect 1230 61019 1286 61075
rect 1354 61019 1410 61075
rect 1478 61019 1534 61075
rect 1602 61019 1658 61075
rect 1726 61019 1782 61075
rect 1850 61019 1906 61075
rect 114 60895 170 60951
rect 238 60895 294 60951
rect 362 60895 418 60951
rect 486 60895 542 60951
rect 610 60895 666 60951
rect 734 60895 790 60951
rect 858 60895 914 60951
rect 982 60895 1038 60951
rect 1106 60895 1162 60951
rect 1230 60895 1286 60951
rect 1354 60895 1410 60951
rect 1478 60895 1534 60951
rect 1602 60895 1658 60951
rect 1726 60895 1782 60951
rect 1850 60895 1906 60951
rect 114 60771 170 60827
rect 238 60771 294 60827
rect 362 60771 418 60827
rect 486 60771 542 60827
rect 610 60771 666 60827
rect 734 60771 790 60827
rect 858 60771 914 60827
rect 982 60771 1038 60827
rect 1106 60771 1162 60827
rect 1230 60771 1286 60827
rect 1354 60771 1410 60827
rect 1478 60771 1534 60827
rect 1602 60771 1658 60827
rect 1726 60771 1782 60827
rect 1850 60771 1906 60827
rect 114 60647 170 60703
rect 238 60647 294 60703
rect 362 60647 418 60703
rect 486 60647 542 60703
rect 610 60647 666 60703
rect 734 60647 790 60703
rect 858 60647 914 60703
rect 982 60647 1038 60703
rect 1106 60647 1162 60703
rect 1230 60647 1286 60703
rect 1354 60647 1410 60703
rect 1478 60647 1534 60703
rect 1602 60647 1658 60703
rect 1726 60647 1782 60703
rect 1850 60647 1906 60703
rect 114 60523 170 60579
rect 238 60523 294 60579
rect 362 60523 418 60579
rect 486 60523 542 60579
rect 610 60523 666 60579
rect 734 60523 790 60579
rect 858 60523 914 60579
rect 982 60523 1038 60579
rect 1106 60523 1162 60579
rect 1230 60523 1286 60579
rect 1354 60523 1410 60579
rect 1478 60523 1534 60579
rect 1602 60523 1658 60579
rect 1726 60523 1782 60579
rect 1850 60523 1906 60579
rect 114 60034 170 60090
rect 238 60034 294 60090
rect 362 60034 418 60090
rect 486 60034 542 60090
rect 610 60034 666 60090
rect 734 60034 790 60090
rect 858 60034 914 60090
rect 982 60034 1038 60090
rect 1106 60034 1162 60090
rect 1230 60034 1286 60090
rect 1354 60034 1410 60090
rect 1478 60034 1534 60090
rect 1602 60034 1658 60090
rect 1726 60034 1782 60090
rect 1850 60034 1906 60090
rect 114 59910 170 59966
rect 238 59910 294 59966
rect 362 59910 418 59966
rect 486 59910 542 59966
rect 610 59910 666 59966
rect 734 59910 790 59966
rect 858 59910 914 59966
rect 982 59910 1038 59966
rect 1106 59910 1162 59966
rect 1230 59910 1286 59966
rect 1354 59910 1410 59966
rect 1478 59910 1534 59966
rect 1602 59910 1658 59966
rect 1726 59910 1782 59966
rect 1850 59910 1906 59966
rect 114 59786 170 59842
rect 238 59786 294 59842
rect 362 59786 418 59842
rect 486 59786 542 59842
rect 610 59786 666 59842
rect 734 59786 790 59842
rect 858 59786 914 59842
rect 982 59786 1038 59842
rect 1106 59786 1162 59842
rect 1230 59786 1286 59842
rect 1354 59786 1410 59842
rect 1478 59786 1534 59842
rect 1602 59786 1658 59842
rect 1726 59786 1782 59842
rect 1850 59786 1906 59842
rect 114 59662 170 59718
rect 238 59662 294 59718
rect 362 59662 418 59718
rect 486 59662 542 59718
rect 610 59662 666 59718
rect 734 59662 790 59718
rect 858 59662 914 59718
rect 982 59662 1038 59718
rect 1106 59662 1162 59718
rect 1230 59662 1286 59718
rect 1354 59662 1410 59718
rect 1478 59662 1534 59718
rect 1602 59662 1658 59718
rect 1726 59662 1782 59718
rect 1850 59662 1906 59718
rect 114 59538 170 59594
rect 238 59538 294 59594
rect 362 59538 418 59594
rect 486 59538 542 59594
rect 610 59538 666 59594
rect 734 59538 790 59594
rect 858 59538 914 59594
rect 982 59538 1038 59594
rect 1106 59538 1162 59594
rect 1230 59538 1286 59594
rect 1354 59538 1410 59594
rect 1478 59538 1534 59594
rect 1602 59538 1658 59594
rect 1726 59538 1782 59594
rect 1850 59538 1906 59594
rect 114 59414 170 59470
rect 238 59414 294 59470
rect 362 59414 418 59470
rect 486 59414 542 59470
rect 610 59414 666 59470
rect 734 59414 790 59470
rect 858 59414 914 59470
rect 982 59414 1038 59470
rect 1106 59414 1162 59470
rect 1230 59414 1286 59470
rect 1354 59414 1410 59470
rect 1478 59414 1534 59470
rect 1602 59414 1658 59470
rect 1726 59414 1782 59470
rect 1850 59414 1906 59470
rect 114 59290 170 59346
rect 238 59290 294 59346
rect 362 59290 418 59346
rect 486 59290 542 59346
rect 610 59290 666 59346
rect 734 59290 790 59346
rect 858 59290 914 59346
rect 982 59290 1038 59346
rect 1106 59290 1162 59346
rect 1230 59290 1286 59346
rect 1354 59290 1410 59346
rect 1478 59290 1534 59346
rect 1602 59290 1658 59346
rect 1726 59290 1782 59346
rect 1850 59290 1906 59346
rect 114 59166 170 59222
rect 238 59166 294 59222
rect 362 59166 418 59222
rect 486 59166 542 59222
rect 610 59166 666 59222
rect 734 59166 790 59222
rect 858 59166 914 59222
rect 982 59166 1038 59222
rect 1106 59166 1162 59222
rect 1230 59166 1286 59222
rect 1354 59166 1410 59222
rect 1478 59166 1534 59222
rect 1602 59166 1658 59222
rect 1726 59166 1782 59222
rect 1850 59166 1906 59222
rect 114 59042 170 59098
rect 238 59042 294 59098
rect 362 59042 418 59098
rect 486 59042 542 59098
rect 610 59042 666 59098
rect 734 59042 790 59098
rect 858 59042 914 59098
rect 982 59042 1038 59098
rect 1106 59042 1162 59098
rect 1230 59042 1286 59098
rect 1354 59042 1410 59098
rect 1478 59042 1534 59098
rect 1602 59042 1658 59098
rect 1726 59042 1782 59098
rect 1850 59042 1906 59098
rect 114 58918 170 58974
rect 238 58918 294 58974
rect 362 58918 418 58974
rect 486 58918 542 58974
rect 610 58918 666 58974
rect 734 58918 790 58974
rect 858 58918 914 58974
rect 982 58918 1038 58974
rect 1106 58918 1162 58974
rect 1230 58918 1286 58974
rect 1354 58918 1410 58974
rect 1478 58918 1534 58974
rect 1602 58918 1658 58974
rect 1726 58918 1782 58974
rect 1850 58918 1906 58974
rect 114 58429 170 58485
rect 238 58429 294 58485
rect 362 58429 418 58485
rect 486 58429 542 58485
rect 610 58429 666 58485
rect 734 58429 790 58485
rect 858 58429 914 58485
rect 982 58429 1038 58485
rect 1106 58429 1162 58485
rect 1230 58429 1286 58485
rect 1354 58429 1410 58485
rect 1478 58429 1534 58485
rect 1602 58429 1658 58485
rect 1726 58429 1782 58485
rect 1850 58429 1906 58485
rect 114 58305 170 58361
rect 238 58305 294 58361
rect 362 58305 418 58361
rect 486 58305 542 58361
rect 610 58305 666 58361
rect 734 58305 790 58361
rect 858 58305 914 58361
rect 982 58305 1038 58361
rect 1106 58305 1162 58361
rect 1230 58305 1286 58361
rect 1354 58305 1410 58361
rect 1478 58305 1534 58361
rect 1602 58305 1658 58361
rect 1726 58305 1782 58361
rect 1850 58305 1906 58361
rect 114 58181 170 58237
rect 238 58181 294 58237
rect 362 58181 418 58237
rect 486 58181 542 58237
rect 610 58181 666 58237
rect 734 58181 790 58237
rect 858 58181 914 58237
rect 982 58181 1038 58237
rect 1106 58181 1162 58237
rect 1230 58181 1286 58237
rect 1354 58181 1410 58237
rect 1478 58181 1534 58237
rect 1602 58181 1658 58237
rect 1726 58181 1782 58237
rect 1850 58181 1906 58237
rect 114 58057 170 58113
rect 238 58057 294 58113
rect 362 58057 418 58113
rect 486 58057 542 58113
rect 610 58057 666 58113
rect 734 58057 790 58113
rect 858 58057 914 58113
rect 982 58057 1038 58113
rect 1106 58057 1162 58113
rect 1230 58057 1286 58113
rect 1354 58057 1410 58113
rect 1478 58057 1534 58113
rect 1602 58057 1658 58113
rect 1726 58057 1782 58113
rect 1850 58057 1906 58113
rect 114 57933 170 57989
rect 238 57933 294 57989
rect 362 57933 418 57989
rect 486 57933 542 57989
rect 610 57933 666 57989
rect 734 57933 790 57989
rect 858 57933 914 57989
rect 982 57933 1038 57989
rect 1106 57933 1162 57989
rect 1230 57933 1286 57989
rect 1354 57933 1410 57989
rect 1478 57933 1534 57989
rect 1602 57933 1658 57989
rect 1726 57933 1782 57989
rect 1850 57933 1906 57989
rect 114 57809 170 57865
rect 238 57809 294 57865
rect 362 57809 418 57865
rect 486 57809 542 57865
rect 610 57809 666 57865
rect 734 57809 790 57865
rect 858 57809 914 57865
rect 982 57809 1038 57865
rect 1106 57809 1162 57865
rect 1230 57809 1286 57865
rect 1354 57809 1410 57865
rect 1478 57809 1534 57865
rect 1602 57809 1658 57865
rect 1726 57809 1782 57865
rect 1850 57809 1906 57865
rect 114 57685 170 57741
rect 238 57685 294 57741
rect 362 57685 418 57741
rect 486 57685 542 57741
rect 610 57685 666 57741
rect 734 57685 790 57741
rect 858 57685 914 57741
rect 982 57685 1038 57741
rect 1106 57685 1162 57741
rect 1230 57685 1286 57741
rect 1354 57685 1410 57741
rect 1478 57685 1534 57741
rect 1602 57685 1658 57741
rect 1726 57685 1782 57741
rect 1850 57685 1906 57741
rect 114 57561 170 57617
rect 238 57561 294 57617
rect 362 57561 418 57617
rect 486 57561 542 57617
rect 610 57561 666 57617
rect 734 57561 790 57617
rect 858 57561 914 57617
rect 982 57561 1038 57617
rect 1106 57561 1162 57617
rect 1230 57561 1286 57617
rect 1354 57561 1410 57617
rect 1478 57561 1534 57617
rect 1602 57561 1658 57617
rect 1726 57561 1782 57617
rect 1850 57561 1906 57617
rect 114 57437 170 57493
rect 238 57437 294 57493
rect 362 57437 418 57493
rect 486 57437 542 57493
rect 610 57437 666 57493
rect 734 57437 790 57493
rect 858 57437 914 57493
rect 982 57437 1038 57493
rect 1106 57437 1162 57493
rect 1230 57437 1286 57493
rect 1354 57437 1410 57493
rect 1478 57437 1534 57493
rect 1602 57437 1658 57493
rect 1726 57437 1782 57493
rect 1850 57437 1906 57493
rect 114 57313 170 57369
rect 238 57313 294 57369
rect 362 57313 418 57369
rect 486 57313 542 57369
rect 610 57313 666 57369
rect 734 57313 790 57369
rect 858 57313 914 57369
rect 982 57313 1038 57369
rect 1106 57313 1162 57369
rect 1230 57313 1286 57369
rect 1354 57313 1410 57369
rect 1478 57313 1534 57369
rect 1602 57313 1658 57369
rect 1726 57313 1782 57369
rect 1850 57313 1906 57369
rect 114 56833 170 56889
rect 238 56833 294 56889
rect 362 56833 418 56889
rect 486 56833 542 56889
rect 610 56833 666 56889
rect 734 56833 790 56889
rect 858 56833 914 56889
rect 982 56833 1038 56889
rect 1106 56833 1162 56889
rect 1230 56833 1286 56889
rect 1354 56833 1410 56889
rect 1478 56833 1534 56889
rect 1602 56833 1658 56889
rect 1726 56833 1782 56889
rect 1850 56833 1906 56889
rect 114 56709 170 56765
rect 238 56709 294 56765
rect 362 56709 418 56765
rect 486 56709 542 56765
rect 610 56709 666 56765
rect 734 56709 790 56765
rect 858 56709 914 56765
rect 982 56709 1038 56765
rect 1106 56709 1162 56765
rect 1230 56709 1286 56765
rect 1354 56709 1410 56765
rect 1478 56709 1534 56765
rect 1602 56709 1658 56765
rect 1726 56709 1782 56765
rect 1850 56709 1906 56765
rect 114 56585 170 56641
rect 238 56585 294 56641
rect 362 56585 418 56641
rect 486 56585 542 56641
rect 610 56585 666 56641
rect 734 56585 790 56641
rect 858 56585 914 56641
rect 982 56585 1038 56641
rect 1106 56585 1162 56641
rect 1230 56585 1286 56641
rect 1354 56585 1410 56641
rect 1478 56585 1534 56641
rect 1602 56585 1658 56641
rect 1726 56585 1782 56641
rect 1850 56585 1906 56641
rect 114 56461 170 56517
rect 238 56461 294 56517
rect 362 56461 418 56517
rect 486 56461 542 56517
rect 610 56461 666 56517
rect 734 56461 790 56517
rect 858 56461 914 56517
rect 982 56461 1038 56517
rect 1106 56461 1162 56517
rect 1230 56461 1286 56517
rect 1354 56461 1410 56517
rect 1478 56461 1534 56517
rect 1602 56461 1658 56517
rect 1726 56461 1782 56517
rect 1850 56461 1906 56517
rect 114 56337 170 56393
rect 238 56337 294 56393
rect 362 56337 418 56393
rect 486 56337 542 56393
rect 610 56337 666 56393
rect 734 56337 790 56393
rect 858 56337 914 56393
rect 982 56337 1038 56393
rect 1106 56337 1162 56393
rect 1230 56337 1286 56393
rect 1354 56337 1410 56393
rect 1478 56337 1534 56393
rect 1602 56337 1658 56393
rect 1726 56337 1782 56393
rect 1850 56337 1906 56393
rect 114 56213 170 56269
rect 238 56213 294 56269
rect 362 56213 418 56269
rect 486 56213 542 56269
rect 610 56213 666 56269
rect 734 56213 790 56269
rect 858 56213 914 56269
rect 982 56213 1038 56269
rect 1106 56213 1162 56269
rect 1230 56213 1286 56269
rect 1354 56213 1410 56269
rect 1478 56213 1534 56269
rect 1602 56213 1658 56269
rect 1726 56213 1782 56269
rect 1850 56213 1906 56269
rect 114 56089 170 56145
rect 238 56089 294 56145
rect 362 56089 418 56145
rect 486 56089 542 56145
rect 610 56089 666 56145
rect 734 56089 790 56145
rect 858 56089 914 56145
rect 982 56089 1038 56145
rect 1106 56089 1162 56145
rect 1230 56089 1286 56145
rect 1354 56089 1410 56145
rect 1478 56089 1534 56145
rect 1602 56089 1658 56145
rect 1726 56089 1782 56145
rect 1850 56089 1906 56145
rect 114 55965 170 56021
rect 238 55965 294 56021
rect 362 55965 418 56021
rect 486 55965 542 56021
rect 610 55965 666 56021
rect 734 55965 790 56021
rect 858 55965 914 56021
rect 982 55965 1038 56021
rect 1106 55965 1162 56021
rect 1230 55965 1286 56021
rect 1354 55965 1410 56021
rect 1478 55965 1534 56021
rect 1602 55965 1658 56021
rect 1726 55965 1782 56021
rect 1850 55965 1906 56021
rect 114 55841 170 55897
rect 238 55841 294 55897
rect 362 55841 418 55897
rect 486 55841 542 55897
rect 610 55841 666 55897
rect 734 55841 790 55897
rect 858 55841 914 55897
rect 982 55841 1038 55897
rect 1106 55841 1162 55897
rect 1230 55841 1286 55897
rect 1354 55841 1410 55897
rect 1478 55841 1534 55897
rect 1602 55841 1658 55897
rect 1726 55841 1782 55897
rect 1850 55841 1906 55897
rect 114 55717 170 55773
rect 238 55717 294 55773
rect 362 55717 418 55773
rect 486 55717 542 55773
rect 610 55717 666 55773
rect 734 55717 790 55773
rect 858 55717 914 55773
rect 982 55717 1038 55773
rect 1106 55717 1162 55773
rect 1230 55717 1286 55773
rect 1354 55717 1410 55773
rect 1478 55717 1534 55773
rect 1602 55717 1658 55773
rect 1726 55717 1782 55773
rect 1850 55717 1906 55773
rect 114 55224 170 55280
rect 238 55224 294 55280
rect 362 55224 418 55280
rect 486 55224 542 55280
rect 610 55224 666 55280
rect 734 55224 790 55280
rect 858 55224 914 55280
rect 982 55224 1038 55280
rect 1106 55224 1162 55280
rect 1230 55224 1286 55280
rect 1354 55224 1410 55280
rect 1478 55224 1534 55280
rect 1602 55224 1658 55280
rect 1726 55224 1782 55280
rect 1850 55224 1906 55280
rect 114 55100 170 55156
rect 238 55100 294 55156
rect 362 55100 418 55156
rect 486 55100 542 55156
rect 610 55100 666 55156
rect 734 55100 790 55156
rect 858 55100 914 55156
rect 982 55100 1038 55156
rect 1106 55100 1162 55156
rect 1230 55100 1286 55156
rect 1354 55100 1410 55156
rect 1478 55100 1534 55156
rect 1602 55100 1658 55156
rect 1726 55100 1782 55156
rect 1850 55100 1906 55156
rect 114 54976 170 55032
rect 238 54976 294 55032
rect 362 54976 418 55032
rect 486 54976 542 55032
rect 610 54976 666 55032
rect 734 54976 790 55032
rect 858 54976 914 55032
rect 982 54976 1038 55032
rect 1106 54976 1162 55032
rect 1230 54976 1286 55032
rect 1354 54976 1410 55032
rect 1478 54976 1534 55032
rect 1602 54976 1658 55032
rect 1726 54976 1782 55032
rect 1850 54976 1906 55032
rect 114 54852 170 54908
rect 238 54852 294 54908
rect 362 54852 418 54908
rect 486 54852 542 54908
rect 610 54852 666 54908
rect 734 54852 790 54908
rect 858 54852 914 54908
rect 982 54852 1038 54908
rect 1106 54852 1162 54908
rect 1230 54852 1286 54908
rect 1354 54852 1410 54908
rect 1478 54852 1534 54908
rect 1602 54852 1658 54908
rect 1726 54852 1782 54908
rect 1850 54852 1906 54908
rect 114 54728 170 54784
rect 238 54728 294 54784
rect 362 54728 418 54784
rect 486 54728 542 54784
rect 610 54728 666 54784
rect 734 54728 790 54784
rect 858 54728 914 54784
rect 982 54728 1038 54784
rect 1106 54728 1162 54784
rect 1230 54728 1286 54784
rect 1354 54728 1410 54784
rect 1478 54728 1534 54784
rect 1602 54728 1658 54784
rect 1726 54728 1782 54784
rect 1850 54728 1906 54784
rect 114 54604 170 54660
rect 238 54604 294 54660
rect 362 54604 418 54660
rect 486 54604 542 54660
rect 610 54604 666 54660
rect 734 54604 790 54660
rect 858 54604 914 54660
rect 982 54604 1038 54660
rect 1106 54604 1162 54660
rect 1230 54604 1286 54660
rect 1354 54604 1410 54660
rect 1478 54604 1534 54660
rect 1602 54604 1658 54660
rect 1726 54604 1782 54660
rect 1850 54604 1906 54660
rect 114 54480 170 54536
rect 238 54480 294 54536
rect 362 54480 418 54536
rect 486 54480 542 54536
rect 610 54480 666 54536
rect 734 54480 790 54536
rect 858 54480 914 54536
rect 982 54480 1038 54536
rect 1106 54480 1162 54536
rect 1230 54480 1286 54536
rect 1354 54480 1410 54536
rect 1478 54480 1534 54536
rect 1602 54480 1658 54536
rect 1726 54480 1782 54536
rect 1850 54480 1906 54536
rect 114 54356 170 54412
rect 238 54356 294 54412
rect 362 54356 418 54412
rect 486 54356 542 54412
rect 610 54356 666 54412
rect 734 54356 790 54412
rect 858 54356 914 54412
rect 982 54356 1038 54412
rect 1106 54356 1162 54412
rect 1230 54356 1286 54412
rect 1354 54356 1410 54412
rect 1478 54356 1534 54412
rect 1602 54356 1658 54412
rect 1726 54356 1782 54412
rect 1850 54356 1906 54412
rect 114 54232 170 54288
rect 238 54232 294 54288
rect 362 54232 418 54288
rect 486 54232 542 54288
rect 610 54232 666 54288
rect 734 54232 790 54288
rect 858 54232 914 54288
rect 982 54232 1038 54288
rect 1106 54232 1162 54288
rect 1230 54232 1286 54288
rect 1354 54232 1410 54288
rect 1478 54232 1534 54288
rect 1602 54232 1658 54288
rect 1726 54232 1782 54288
rect 1850 54232 1906 54288
rect 114 54108 170 54164
rect 238 54108 294 54164
rect 362 54108 418 54164
rect 486 54108 542 54164
rect 610 54108 666 54164
rect 734 54108 790 54164
rect 858 54108 914 54164
rect 982 54108 1038 54164
rect 1106 54108 1162 54164
rect 1230 54108 1286 54164
rect 1354 54108 1410 54164
rect 1478 54108 1534 54164
rect 1602 54108 1658 54164
rect 1726 54108 1782 54164
rect 1850 54108 1906 54164
rect 114 53651 170 53707
rect 238 53651 294 53707
rect 362 53651 418 53707
rect 486 53651 542 53707
rect 610 53651 666 53707
rect 734 53651 790 53707
rect 858 53651 914 53707
rect 982 53651 1038 53707
rect 1106 53651 1162 53707
rect 1230 53651 1286 53707
rect 1354 53651 1410 53707
rect 1478 53651 1534 53707
rect 1602 53651 1658 53707
rect 1726 53651 1782 53707
rect 1850 53651 1906 53707
rect 114 53527 170 53583
rect 238 53527 294 53583
rect 362 53527 418 53583
rect 486 53527 542 53583
rect 610 53527 666 53583
rect 734 53527 790 53583
rect 858 53527 914 53583
rect 982 53527 1038 53583
rect 1106 53527 1162 53583
rect 1230 53527 1286 53583
rect 1354 53527 1410 53583
rect 1478 53527 1534 53583
rect 1602 53527 1658 53583
rect 1726 53527 1782 53583
rect 1850 53527 1906 53583
rect 114 53403 170 53459
rect 238 53403 294 53459
rect 362 53403 418 53459
rect 486 53403 542 53459
rect 610 53403 666 53459
rect 734 53403 790 53459
rect 858 53403 914 53459
rect 982 53403 1038 53459
rect 1106 53403 1162 53459
rect 1230 53403 1286 53459
rect 1354 53403 1410 53459
rect 1478 53403 1534 53459
rect 1602 53403 1658 53459
rect 1726 53403 1782 53459
rect 1850 53403 1906 53459
rect 114 53279 170 53335
rect 238 53279 294 53335
rect 362 53279 418 53335
rect 486 53279 542 53335
rect 610 53279 666 53335
rect 734 53279 790 53335
rect 858 53279 914 53335
rect 982 53279 1038 53335
rect 1106 53279 1162 53335
rect 1230 53279 1286 53335
rect 1354 53279 1410 53335
rect 1478 53279 1534 53335
rect 1602 53279 1658 53335
rect 1726 53279 1782 53335
rect 1850 53279 1906 53335
rect 114 53155 170 53211
rect 238 53155 294 53211
rect 362 53155 418 53211
rect 486 53155 542 53211
rect 610 53155 666 53211
rect 734 53155 790 53211
rect 858 53155 914 53211
rect 982 53155 1038 53211
rect 1106 53155 1162 53211
rect 1230 53155 1286 53211
rect 1354 53155 1410 53211
rect 1478 53155 1534 53211
rect 1602 53155 1658 53211
rect 1726 53155 1782 53211
rect 1850 53155 1906 53211
rect 114 53031 170 53087
rect 238 53031 294 53087
rect 362 53031 418 53087
rect 486 53031 542 53087
rect 610 53031 666 53087
rect 734 53031 790 53087
rect 858 53031 914 53087
rect 982 53031 1038 53087
rect 1106 53031 1162 53087
rect 1230 53031 1286 53087
rect 1354 53031 1410 53087
rect 1478 53031 1534 53087
rect 1602 53031 1658 53087
rect 1726 53031 1782 53087
rect 1850 53031 1906 53087
rect 114 52907 170 52963
rect 238 52907 294 52963
rect 362 52907 418 52963
rect 486 52907 542 52963
rect 610 52907 666 52963
rect 734 52907 790 52963
rect 858 52907 914 52963
rect 982 52907 1038 52963
rect 1106 52907 1162 52963
rect 1230 52907 1286 52963
rect 1354 52907 1410 52963
rect 1478 52907 1534 52963
rect 1602 52907 1658 52963
rect 1726 52907 1782 52963
rect 1850 52907 1906 52963
rect 114 52783 170 52839
rect 238 52783 294 52839
rect 362 52783 418 52839
rect 486 52783 542 52839
rect 610 52783 666 52839
rect 734 52783 790 52839
rect 858 52783 914 52839
rect 982 52783 1038 52839
rect 1106 52783 1162 52839
rect 1230 52783 1286 52839
rect 1354 52783 1410 52839
rect 1478 52783 1534 52839
rect 1602 52783 1658 52839
rect 1726 52783 1782 52839
rect 1850 52783 1906 52839
rect 114 52659 170 52715
rect 238 52659 294 52715
rect 362 52659 418 52715
rect 486 52659 542 52715
rect 610 52659 666 52715
rect 734 52659 790 52715
rect 858 52659 914 52715
rect 982 52659 1038 52715
rect 1106 52659 1162 52715
rect 1230 52659 1286 52715
rect 1354 52659 1410 52715
rect 1478 52659 1534 52715
rect 1602 52659 1658 52715
rect 1726 52659 1782 52715
rect 1850 52659 1906 52715
rect 114 52535 170 52591
rect 238 52535 294 52591
rect 362 52535 418 52591
rect 486 52535 542 52591
rect 610 52535 666 52591
rect 734 52535 790 52591
rect 858 52535 914 52591
rect 982 52535 1038 52591
rect 1106 52535 1162 52591
rect 1230 52535 1286 52591
rect 1354 52535 1410 52591
rect 1478 52535 1534 52591
rect 1602 52535 1658 52591
rect 1726 52535 1782 52591
rect 1850 52535 1906 52591
rect 114 52044 170 52100
rect 238 52044 294 52100
rect 362 52044 418 52100
rect 486 52044 542 52100
rect 610 52044 666 52100
rect 734 52044 790 52100
rect 858 52044 914 52100
rect 982 52044 1038 52100
rect 1106 52044 1162 52100
rect 1230 52044 1286 52100
rect 1354 52044 1410 52100
rect 1478 52044 1534 52100
rect 1602 52044 1658 52100
rect 1726 52044 1782 52100
rect 1850 52044 1906 52100
rect 114 51920 170 51976
rect 238 51920 294 51976
rect 362 51920 418 51976
rect 486 51920 542 51976
rect 610 51920 666 51976
rect 734 51920 790 51976
rect 858 51920 914 51976
rect 982 51920 1038 51976
rect 1106 51920 1162 51976
rect 1230 51920 1286 51976
rect 1354 51920 1410 51976
rect 1478 51920 1534 51976
rect 1602 51920 1658 51976
rect 1726 51920 1782 51976
rect 1850 51920 1906 51976
rect 114 51796 170 51852
rect 238 51796 294 51852
rect 362 51796 418 51852
rect 486 51796 542 51852
rect 610 51796 666 51852
rect 734 51796 790 51852
rect 858 51796 914 51852
rect 982 51796 1038 51852
rect 1106 51796 1162 51852
rect 1230 51796 1286 51852
rect 1354 51796 1410 51852
rect 1478 51796 1534 51852
rect 1602 51796 1658 51852
rect 1726 51796 1782 51852
rect 1850 51796 1906 51852
rect 114 51672 170 51728
rect 238 51672 294 51728
rect 362 51672 418 51728
rect 486 51672 542 51728
rect 610 51672 666 51728
rect 734 51672 790 51728
rect 858 51672 914 51728
rect 982 51672 1038 51728
rect 1106 51672 1162 51728
rect 1230 51672 1286 51728
rect 1354 51672 1410 51728
rect 1478 51672 1534 51728
rect 1602 51672 1658 51728
rect 1726 51672 1782 51728
rect 1850 51672 1906 51728
rect 114 51548 170 51604
rect 238 51548 294 51604
rect 362 51548 418 51604
rect 486 51548 542 51604
rect 610 51548 666 51604
rect 734 51548 790 51604
rect 858 51548 914 51604
rect 982 51548 1038 51604
rect 1106 51548 1162 51604
rect 1230 51548 1286 51604
rect 1354 51548 1410 51604
rect 1478 51548 1534 51604
rect 1602 51548 1658 51604
rect 1726 51548 1782 51604
rect 1850 51548 1906 51604
rect 114 51424 170 51480
rect 238 51424 294 51480
rect 362 51424 418 51480
rect 486 51424 542 51480
rect 610 51424 666 51480
rect 734 51424 790 51480
rect 858 51424 914 51480
rect 982 51424 1038 51480
rect 1106 51424 1162 51480
rect 1230 51424 1286 51480
rect 1354 51424 1410 51480
rect 1478 51424 1534 51480
rect 1602 51424 1658 51480
rect 1726 51424 1782 51480
rect 1850 51424 1906 51480
rect 114 51300 170 51356
rect 238 51300 294 51356
rect 362 51300 418 51356
rect 486 51300 542 51356
rect 610 51300 666 51356
rect 734 51300 790 51356
rect 858 51300 914 51356
rect 982 51300 1038 51356
rect 1106 51300 1162 51356
rect 1230 51300 1286 51356
rect 1354 51300 1410 51356
rect 1478 51300 1534 51356
rect 1602 51300 1658 51356
rect 1726 51300 1782 51356
rect 1850 51300 1906 51356
rect 114 51176 170 51232
rect 238 51176 294 51232
rect 362 51176 418 51232
rect 486 51176 542 51232
rect 610 51176 666 51232
rect 734 51176 790 51232
rect 858 51176 914 51232
rect 982 51176 1038 51232
rect 1106 51176 1162 51232
rect 1230 51176 1286 51232
rect 1354 51176 1410 51232
rect 1478 51176 1534 51232
rect 1602 51176 1658 51232
rect 1726 51176 1782 51232
rect 1850 51176 1906 51232
rect 114 51052 170 51108
rect 238 51052 294 51108
rect 362 51052 418 51108
rect 486 51052 542 51108
rect 610 51052 666 51108
rect 734 51052 790 51108
rect 858 51052 914 51108
rect 982 51052 1038 51108
rect 1106 51052 1162 51108
rect 1230 51052 1286 51108
rect 1354 51052 1410 51108
rect 1478 51052 1534 51108
rect 1602 51052 1658 51108
rect 1726 51052 1782 51108
rect 1850 51052 1906 51108
rect 114 50928 170 50984
rect 238 50928 294 50984
rect 362 50928 418 50984
rect 486 50928 542 50984
rect 610 50928 666 50984
rect 734 50928 790 50984
rect 858 50928 914 50984
rect 982 50928 1038 50984
rect 1106 50928 1162 50984
rect 1230 50928 1286 50984
rect 1354 50928 1410 50984
rect 1478 50928 1534 50984
rect 1602 50928 1658 50984
rect 1726 50928 1782 50984
rect 1850 50928 1906 50984
rect 114 50424 170 50480
rect 238 50424 294 50480
rect 362 50424 418 50480
rect 486 50424 542 50480
rect 610 50424 666 50480
rect 734 50424 790 50480
rect 858 50424 914 50480
rect 982 50424 1038 50480
rect 1106 50424 1162 50480
rect 1230 50424 1286 50480
rect 1354 50424 1410 50480
rect 1478 50424 1534 50480
rect 1602 50424 1658 50480
rect 1726 50424 1782 50480
rect 1850 50424 1906 50480
rect 114 50300 170 50356
rect 238 50300 294 50356
rect 362 50300 418 50356
rect 486 50300 542 50356
rect 610 50300 666 50356
rect 734 50300 790 50356
rect 858 50300 914 50356
rect 982 50300 1038 50356
rect 1106 50300 1162 50356
rect 1230 50300 1286 50356
rect 1354 50300 1410 50356
rect 1478 50300 1534 50356
rect 1602 50300 1658 50356
rect 1726 50300 1782 50356
rect 1850 50300 1906 50356
rect 114 50176 170 50232
rect 238 50176 294 50232
rect 362 50176 418 50232
rect 486 50176 542 50232
rect 610 50176 666 50232
rect 734 50176 790 50232
rect 858 50176 914 50232
rect 982 50176 1038 50232
rect 1106 50176 1162 50232
rect 1230 50176 1286 50232
rect 1354 50176 1410 50232
rect 1478 50176 1534 50232
rect 1602 50176 1658 50232
rect 1726 50176 1782 50232
rect 1850 50176 1906 50232
rect 114 50052 170 50108
rect 238 50052 294 50108
rect 362 50052 418 50108
rect 486 50052 542 50108
rect 610 50052 666 50108
rect 734 50052 790 50108
rect 858 50052 914 50108
rect 982 50052 1038 50108
rect 1106 50052 1162 50108
rect 1230 50052 1286 50108
rect 1354 50052 1410 50108
rect 1478 50052 1534 50108
rect 1602 50052 1658 50108
rect 1726 50052 1782 50108
rect 1850 50052 1906 50108
rect 114 49928 170 49984
rect 238 49928 294 49984
rect 362 49928 418 49984
rect 486 49928 542 49984
rect 610 49928 666 49984
rect 734 49928 790 49984
rect 858 49928 914 49984
rect 982 49928 1038 49984
rect 1106 49928 1162 49984
rect 1230 49928 1286 49984
rect 1354 49928 1410 49984
rect 1478 49928 1534 49984
rect 1602 49928 1658 49984
rect 1726 49928 1782 49984
rect 1850 49928 1906 49984
rect 114 49804 170 49860
rect 238 49804 294 49860
rect 362 49804 418 49860
rect 486 49804 542 49860
rect 610 49804 666 49860
rect 734 49804 790 49860
rect 858 49804 914 49860
rect 982 49804 1038 49860
rect 1106 49804 1162 49860
rect 1230 49804 1286 49860
rect 1354 49804 1410 49860
rect 1478 49804 1534 49860
rect 1602 49804 1658 49860
rect 1726 49804 1782 49860
rect 1850 49804 1906 49860
rect 114 49680 170 49736
rect 238 49680 294 49736
rect 362 49680 418 49736
rect 486 49680 542 49736
rect 610 49680 666 49736
rect 734 49680 790 49736
rect 858 49680 914 49736
rect 982 49680 1038 49736
rect 1106 49680 1162 49736
rect 1230 49680 1286 49736
rect 1354 49680 1410 49736
rect 1478 49680 1534 49736
rect 1602 49680 1658 49736
rect 1726 49680 1782 49736
rect 1850 49680 1906 49736
rect 114 49556 170 49612
rect 238 49556 294 49612
rect 362 49556 418 49612
rect 486 49556 542 49612
rect 610 49556 666 49612
rect 734 49556 790 49612
rect 858 49556 914 49612
rect 982 49556 1038 49612
rect 1106 49556 1162 49612
rect 1230 49556 1286 49612
rect 1354 49556 1410 49612
rect 1478 49556 1534 49612
rect 1602 49556 1658 49612
rect 1726 49556 1782 49612
rect 1850 49556 1906 49612
rect 114 49432 170 49488
rect 238 49432 294 49488
rect 362 49432 418 49488
rect 486 49432 542 49488
rect 610 49432 666 49488
rect 734 49432 790 49488
rect 858 49432 914 49488
rect 982 49432 1038 49488
rect 1106 49432 1162 49488
rect 1230 49432 1286 49488
rect 1354 49432 1410 49488
rect 1478 49432 1534 49488
rect 1602 49432 1658 49488
rect 1726 49432 1782 49488
rect 1850 49432 1906 49488
rect 114 49308 170 49364
rect 238 49308 294 49364
rect 362 49308 418 49364
rect 486 49308 542 49364
rect 610 49308 666 49364
rect 734 49308 790 49364
rect 858 49308 914 49364
rect 982 49308 1038 49364
rect 1106 49308 1162 49364
rect 1230 49308 1286 49364
rect 1354 49308 1410 49364
rect 1478 49308 1534 49364
rect 1602 49308 1658 49364
rect 1726 49308 1782 49364
rect 1850 49308 1906 49364
rect 114 48785 170 48841
rect 238 48785 294 48841
rect 362 48785 418 48841
rect 486 48785 542 48841
rect 610 48785 666 48841
rect 734 48785 790 48841
rect 858 48785 914 48841
rect 982 48785 1038 48841
rect 1106 48785 1162 48841
rect 1230 48785 1286 48841
rect 1354 48785 1410 48841
rect 1478 48785 1534 48841
rect 1602 48785 1658 48841
rect 1726 48785 1782 48841
rect 1850 48785 1906 48841
rect 114 48661 170 48717
rect 238 48661 294 48717
rect 362 48661 418 48717
rect 486 48661 542 48717
rect 610 48661 666 48717
rect 734 48661 790 48717
rect 858 48661 914 48717
rect 982 48661 1038 48717
rect 1106 48661 1162 48717
rect 1230 48661 1286 48717
rect 1354 48661 1410 48717
rect 1478 48661 1534 48717
rect 1602 48661 1658 48717
rect 1726 48661 1782 48717
rect 1850 48661 1906 48717
rect 114 48537 170 48593
rect 238 48537 294 48593
rect 362 48537 418 48593
rect 486 48537 542 48593
rect 610 48537 666 48593
rect 734 48537 790 48593
rect 858 48537 914 48593
rect 982 48537 1038 48593
rect 1106 48537 1162 48593
rect 1230 48537 1286 48593
rect 1354 48537 1410 48593
rect 1478 48537 1534 48593
rect 1602 48537 1658 48593
rect 1726 48537 1782 48593
rect 1850 48537 1906 48593
rect 114 48413 170 48469
rect 238 48413 294 48469
rect 362 48413 418 48469
rect 486 48413 542 48469
rect 610 48413 666 48469
rect 734 48413 790 48469
rect 858 48413 914 48469
rect 982 48413 1038 48469
rect 1106 48413 1162 48469
rect 1230 48413 1286 48469
rect 1354 48413 1410 48469
rect 1478 48413 1534 48469
rect 1602 48413 1658 48469
rect 1726 48413 1782 48469
rect 1850 48413 1906 48469
rect 114 48289 170 48345
rect 238 48289 294 48345
rect 362 48289 418 48345
rect 486 48289 542 48345
rect 610 48289 666 48345
rect 734 48289 790 48345
rect 858 48289 914 48345
rect 982 48289 1038 48345
rect 1106 48289 1162 48345
rect 1230 48289 1286 48345
rect 1354 48289 1410 48345
rect 1478 48289 1534 48345
rect 1602 48289 1658 48345
rect 1726 48289 1782 48345
rect 1850 48289 1906 48345
rect 114 48165 170 48221
rect 238 48165 294 48221
rect 362 48165 418 48221
rect 486 48165 542 48221
rect 610 48165 666 48221
rect 734 48165 790 48221
rect 858 48165 914 48221
rect 982 48165 1038 48221
rect 1106 48165 1162 48221
rect 1230 48165 1286 48221
rect 1354 48165 1410 48221
rect 1478 48165 1534 48221
rect 1602 48165 1658 48221
rect 1726 48165 1782 48221
rect 1850 48165 1906 48221
rect 114 48041 170 48097
rect 238 48041 294 48097
rect 362 48041 418 48097
rect 486 48041 542 48097
rect 610 48041 666 48097
rect 734 48041 790 48097
rect 858 48041 914 48097
rect 982 48041 1038 48097
rect 1106 48041 1162 48097
rect 1230 48041 1286 48097
rect 1354 48041 1410 48097
rect 1478 48041 1534 48097
rect 1602 48041 1658 48097
rect 1726 48041 1782 48097
rect 1850 48041 1906 48097
rect 114 47917 170 47973
rect 238 47917 294 47973
rect 362 47917 418 47973
rect 486 47917 542 47973
rect 610 47917 666 47973
rect 734 47917 790 47973
rect 858 47917 914 47973
rect 982 47917 1038 47973
rect 1106 47917 1162 47973
rect 1230 47917 1286 47973
rect 1354 47917 1410 47973
rect 1478 47917 1534 47973
rect 1602 47917 1658 47973
rect 1726 47917 1782 47973
rect 1850 47917 1906 47973
rect 114 47793 170 47849
rect 238 47793 294 47849
rect 362 47793 418 47849
rect 486 47793 542 47849
rect 610 47793 666 47849
rect 734 47793 790 47849
rect 858 47793 914 47849
rect 982 47793 1038 47849
rect 1106 47793 1162 47849
rect 1230 47793 1286 47849
rect 1354 47793 1410 47849
rect 1478 47793 1534 47849
rect 1602 47793 1658 47849
rect 1726 47793 1782 47849
rect 1850 47793 1906 47849
rect 114 47669 170 47725
rect 238 47669 294 47725
rect 362 47669 418 47725
rect 486 47669 542 47725
rect 610 47669 666 47725
rect 734 47669 790 47725
rect 858 47669 914 47725
rect 982 47669 1038 47725
rect 1106 47669 1162 47725
rect 1230 47669 1286 47725
rect 1354 47669 1410 47725
rect 1478 47669 1534 47725
rect 1602 47669 1658 47725
rect 1726 47669 1782 47725
rect 1850 47669 1906 47725
rect 114 47545 170 47601
rect 238 47545 294 47601
rect 362 47545 418 47601
rect 486 47545 542 47601
rect 610 47545 666 47601
rect 734 47545 790 47601
rect 858 47545 914 47601
rect 982 47545 1038 47601
rect 1106 47545 1162 47601
rect 1230 47545 1286 47601
rect 1354 47545 1410 47601
rect 1478 47545 1534 47601
rect 1602 47545 1658 47601
rect 1726 47545 1782 47601
rect 1850 47545 1906 47601
rect 114 47421 170 47477
rect 238 47421 294 47477
rect 362 47421 418 47477
rect 486 47421 542 47477
rect 610 47421 666 47477
rect 734 47421 790 47477
rect 858 47421 914 47477
rect 982 47421 1038 47477
rect 1106 47421 1162 47477
rect 1230 47421 1286 47477
rect 1354 47421 1410 47477
rect 1478 47421 1534 47477
rect 1602 47421 1658 47477
rect 1726 47421 1782 47477
rect 1850 47421 1906 47477
rect 114 47297 170 47353
rect 238 47297 294 47353
rect 362 47297 418 47353
rect 486 47297 542 47353
rect 610 47297 666 47353
rect 734 47297 790 47353
rect 858 47297 914 47353
rect 982 47297 1038 47353
rect 1106 47297 1162 47353
rect 1230 47297 1286 47353
rect 1354 47297 1410 47353
rect 1478 47297 1534 47353
rect 1602 47297 1658 47353
rect 1726 47297 1782 47353
rect 1850 47297 1906 47353
rect 114 47173 170 47229
rect 238 47173 294 47229
rect 362 47173 418 47229
rect 486 47173 542 47229
rect 610 47173 666 47229
rect 734 47173 790 47229
rect 858 47173 914 47229
rect 982 47173 1038 47229
rect 1106 47173 1162 47229
rect 1230 47173 1286 47229
rect 1354 47173 1410 47229
rect 1478 47173 1534 47229
rect 1602 47173 1658 47229
rect 1726 47173 1782 47229
rect 1850 47173 1906 47229
rect 114 47049 170 47105
rect 238 47049 294 47105
rect 362 47049 418 47105
rect 486 47049 542 47105
rect 610 47049 666 47105
rect 734 47049 790 47105
rect 858 47049 914 47105
rect 982 47049 1038 47105
rect 1106 47049 1162 47105
rect 1230 47049 1286 47105
rect 1354 47049 1410 47105
rect 1478 47049 1534 47105
rect 1602 47049 1658 47105
rect 1726 47049 1782 47105
rect 1850 47049 1906 47105
rect 114 46925 170 46981
rect 238 46925 294 46981
rect 362 46925 418 46981
rect 486 46925 542 46981
rect 610 46925 666 46981
rect 734 46925 790 46981
rect 858 46925 914 46981
rect 982 46925 1038 46981
rect 1106 46925 1162 46981
rect 1230 46925 1286 46981
rect 1354 46925 1410 46981
rect 1478 46925 1534 46981
rect 1602 46925 1658 46981
rect 1726 46925 1782 46981
rect 1850 46925 1906 46981
rect 114 46801 170 46857
rect 238 46801 294 46857
rect 362 46801 418 46857
rect 486 46801 542 46857
rect 610 46801 666 46857
rect 734 46801 790 46857
rect 858 46801 914 46857
rect 982 46801 1038 46857
rect 1106 46801 1162 46857
rect 1230 46801 1286 46857
rect 1354 46801 1410 46857
rect 1478 46801 1534 46857
rect 1602 46801 1658 46857
rect 1726 46801 1782 46857
rect 1850 46801 1906 46857
rect 114 46677 170 46733
rect 238 46677 294 46733
rect 362 46677 418 46733
rect 486 46677 542 46733
rect 610 46677 666 46733
rect 734 46677 790 46733
rect 858 46677 914 46733
rect 982 46677 1038 46733
rect 1106 46677 1162 46733
rect 1230 46677 1286 46733
rect 1354 46677 1410 46733
rect 1478 46677 1534 46733
rect 1602 46677 1658 46733
rect 1726 46677 1782 46733
rect 1850 46677 1906 46733
rect 114 46553 170 46609
rect 238 46553 294 46609
rect 362 46553 418 46609
rect 486 46553 542 46609
rect 610 46553 666 46609
rect 734 46553 790 46609
rect 858 46553 914 46609
rect 982 46553 1038 46609
rect 1106 46553 1162 46609
rect 1230 46553 1286 46609
rect 1354 46553 1410 46609
rect 1478 46553 1534 46609
rect 1602 46553 1658 46609
rect 1726 46553 1782 46609
rect 1850 46553 1906 46609
rect 114 46429 170 46485
rect 238 46429 294 46485
rect 362 46429 418 46485
rect 486 46429 542 46485
rect 610 46429 666 46485
rect 734 46429 790 46485
rect 858 46429 914 46485
rect 982 46429 1038 46485
rect 1106 46429 1162 46485
rect 1230 46429 1286 46485
rect 1354 46429 1410 46485
rect 1478 46429 1534 46485
rect 1602 46429 1658 46485
rect 1726 46429 1782 46485
rect 1850 46429 1906 46485
rect 114 46305 170 46361
rect 238 46305 294 46361
rect 362 46305 418 46361
rect 486 46305 542 46361
rect 610 46305 666 46361
rect 734 46305 790 46361
rect 858 46305 914 46361
rect 982 46305 1038 46361
rect 1106 46305 1162 46361
rect 1230 46305 1286 46361
rect 1354 46305 1410 46361
rect 1478 46305 1534 46361
rect 1602 46305 1658 46361
rect 1726 46305 1782 46361
rect 1850 46305 1906 46361
rect 114 46181 170 46237
rect 238 46181 294 46237
rect 362 46181 418 46237
rect 486 46181 542 46237
rect 610 46181 666 46237
rect 734 46181 790 46237
rect 858 46181 914 46237
rect 982 46181 1038 46237
rect 1106 46181 1162 46237
rect 1230 46181 1286 46237
rect 1354 46181 1410 46237
rect 1478 46181 1534 46237
rect 1602 46181 1658 46237
rect 1726 46181 1782 46237
rect 1850 46181 1906 46237
rect 114 45596 170 45652
rect 238 45596 294 45652
rect 362 45596 418 45652
rect 486 45596 542 45652
rect 610 45596 666 45652
rect 734 45596 790 45652
rect 858 45596 914 45652
rect 982 45596 1038 45652
rect 1106 45596 1162 45652
rect 1230 45596 1286 45652
rect 1354 45596 1410 45652
rect 1478 45596 1534 45652
rect 1602 45596 1658 45652
rect 1726 45596 1782 45652
rect 1850 45596 1906 45652
rect 114 45472 170 45528
rect 238 45472 294 45528
rect 362 45472 418 45528
rect 486 45472 542 45528
rect 610 45472 666 45528
rect 734 45472 790 45528
rect 858 45472 914 45528
rect 982 45472 1038 45528
rect 1106 45472 1162 45528
rect 1230 45472 1286 45528
rect 1354 45472 1410 45528
rect 1478 45472 1534 45528
rect 1602 45472 1658 45528
rect 1726 45472 1782 45528
rect 1850 45472 1906 45528
rect 114 45348 170 45404
rect 238 45348 294 45404
rect 362 45348 418 45404
rect 486 45348 542 45404
rect 610 45348 666 45404
rect 734 45348 790 45404
rect 858 45348 914 45404
rect 982 45348 1038 45404
rect 1106 45348 1162 45404
rect 1230 45348 1286 45404
rect 1354 45348 1410 45404
rect 1478 45348 1534 45404
rect 1602 45348 1658 45404
rect 1726 45348 1782 45404
rect 1850 45348 1906 45404
rect 114 45224 170 45280
rect 238 45224 294 45280
rect 362 45224 418 45280
rect 486 45224 542 45280
rect 610 45224 666 45280
rect 734 45224 790 45280
rect 858 45224 914 45280
rect 982 45224 1038 45280
rect 1106 45224 1162 45280
rect 1230 45224 1286 45280
rect 1354 45224 1410 45280
rect 1478 45224 1534 45280
rect 1602 45224 1658 45280
rect 1726 45224 1782 45280
rect 1850 45224 1906 45280
rect 114 45100 170 45156
rect 238 45100 294 45156
rect 362 45100 418 45156
rect 486 45100 542 45156
rect 610 45100 666 45156
rect 734 45100 790 45156
rect 858 45100 914 45156
rect 982 45100 1038 45156
rect 1106 45100 1162 45156
rect 1230 45100 1286 45156
rect 1354 45100 1410 45156
rect 1478 45100 1534 45156
rect 1602 45100 1658 45156
rect 1726 45100 1782 45156
rect 1850 45100 1906 45156
rect 114 44976 170 45032
rect 238 44976 294 45032
rect 362 44976 418 45032
rect 486 44976 542 45032
rect 610 44976 666 45032
rect 734 44976 790 45032
rect 858 44976 914 45032
rect 982 44976 1038 45032
rect 1106 44976 1162 45032
rect 1230 44976 1286 45032
rect 1354 44976 1410 45032
rect 1478 44976 1534 45032
rect 1602 44976 1658 45032
rect 1726 44976 1782 45032
rect 1850 44976 1906 45032
rect 114 44852 170 44908
rect 238 44852 294 44908
rect 362 44852 418 44908
rect 486 44852 542 44908
rect 610 44852 666 44908
rect 734 44852 790 44908
rect 858 44852 914 44908
rect 982 44852 1038 44908
rect 1106 44852 1162 44908
rect 1230 44852 1286 44908
rect 1354 44852 1410 44908
rect 1478 44852 1534 44908
rect 1602 44852 1658 44908
rect 1726 44852 1782 44908
rect 1850 44852 1906 44908
rect 114 44728 170 44784
rect 238 44728 294 44784
rect 362 44728 418 44784
rect 486 44728 542 44784
rect 610 44728 666 44784
rect 734 44728 790 44784
rect 858 44728 914 44784
rect 982 44728 1038 44784
rect 1106 44728 1162 44784
rect 1230 44728 1286 44784
rect 1354 44728 1410 44784
rect 1478 44728 1534 44784
rect 1602 44728 1658 44784
rect 1726 44728 1782 44784
rect 1850 44728 1906 44784
rect 114 44604 170 44660
rect 238 44604 294 44660
rect 362 44604 418 44660
rect 486 44604 542 44660
rect 610 44604 666 44660
rect 734 44604 790 44660
rect 858 44604 914 44660
rect 982 44604 1038 44660
rect 1106 44604 1162 44660
rect 1230 44604 1286 44660
rect 1354 44604 1410 44660
rect 1478 44604 1534 44660
rect 1602 44604 1658 44660
rect 1726 44604 1782 44660
rect 1850 44604 1906 44660
rect 114 44480 170 44536
rect 238 44480 294 44536
rect 362 44480 418 44536
rect 486 44480 542 44536
rect 610 44480 666 44536
rect 734 44480 790 44536
rect 858 44480 914 44536
rect 982 44480 1038 44536
rect 1106 44480 1162 44536
rect 1230 44480 1286 44536
rect 1354 44480 1410 44536
rect 1478 44480 1534 44536
rect 1602 44480 1658 44536
rect 1726 44480 1782 44536
rect 1850 44480 1906 44536
rect 114 44356 170 44412
rect 238 44356 294 44412
rect 362 44356 418 44412
rect 486 44356 542 44412
rect 610 44356 666 44412
rect 734 44356 790 44412
rect 858 44356 914 44412
rect 982 44356 1038 44412
rect 1106 44356 1162 44412
rect 1230 44356 1286 44412
rect 1354 44356 1410 44412
rect 1478 44356 1534 44412
rect 1602 44356 1658 44412
rect 1726 44356 1782 44412
rect 1850 44356 1906 44412
rect 114 44232 170 44288
rect 238 44232 294 44288
rect 362 44232 418 44288
rect 486 44232 542 44288
rect 610 44232 666 44288
rect 734 44232 790 44288
rect 858 44232 914 44288
rect 982 44232 1038 44288
rect 1106 44232 1162 44288
rect 1230 44232 1286 44288
rect 1354 44232 1410 44288
rect 1478 44232 1534 44288
rect 1602 44232 1658 44288
rect 1726 44232 1782 44288
rect 1850 44232 1906 44288
rect 114 44108 170 44164
rect 238 44108 294 44164
rect 362 44108 418 44164
rect 486 44108 542 44164
rect 610 44108 666 44164
rect 734 44108 790 44164
rect 858 44108 914 44164
rect 982 44108 1038 44164
rect 1106 44108 1162 44164
rect 1230 44108 1286 44164
rect 1354 44108 1410 44164
rect 1478 44108 1534 44164
rect 1602 44108 1658 44164
rect 1726 44108 1782 44164
rect 1850 44108 1906 44164
rect 114 43984 170 44040
rect 238 43984 294 44040
rect 362 43984 418 44040
rect 486 43984 542 44040
rect 610 43984 666 44040
rect 734 43984 790 44040
rect 858 43984 914 44040
rect 982 43984 1038 44040
rect 1106 43984 1162 44040
rect 1230 43984 1286 44040
rect 1354 43984 1410 44040
rect 1478 43984 1534 44040
rect 1602 43984 1658 44040
rect 1726 43984 1782 44040
rect 1850 43984 1906 44040
rect 114 43860 170 43916
rect 238 43860 294 43916
rect 362 43860 418 43916
rect 486 43860 542 43916
rect 610 43860 666 43916
rect 734 43860 790 43916
rect 858 43860 914 43916
rect 982 43860 1038 43916
rect 1106 43860 1162 43916
rect 1230 43860 1286 43916
rect 1354 43860 1410 43916
rect 1478 43860 1534 43916
rect 1602 43860 1658 43916
rect 1726 43860 1782 43916
rect 1850 43860 1906 43916
rect 114 43736 170 43792
rect 238 43736 294 43792
rect 362 43736 418 43792
rect 486 43736 542 43792
rect 610 43736 666 43792
rect 734 43736 790 43792
rect 858 43736 914 43792
rect 982 43736 1038 43792
rect 1106 43736 1162 43792
rect 1230 43736 1286 43792
rect 1354 43736 1410 43792
rect 1478 43736 1534 43792
rect 1602 43736 1658 43792
rect 1726 43736 1782 43792
rect 1850 43736 1906 43792
rect 114 43612 170 43668
rect 238 43612 294 43668
rect 362 43612 418 43668
rect 486 43612 542 43668
rect 610 43612 666 43668
rect 734 43612 790 43668
rect 858 43612 914 43668
rect 982 43612 1038 43668
rect 1106 43612 1162 43668
rect 1230 43612 1286 43668
rect 1354 43612 1410 43668
rect 1478 43612 1534 43668
rect 1602 43612 1658 43668
rect 1726 43612 1782 43668
rect 1850 43612 1906 43668
rect 114 43488 170 43544
rect 238 43488 294 43544
rect 362 43488 418 43544
rect 486 43488 542 43544
rect 610 43488 666 43544
rect 734 43488 790 43544
rect 858 43488 914 43544
rect 982 43488 1038 43544
rect 1106 43488 1162 43544
rect 1230 43488 1286 43544
rect 1354 43488 1410 43544
rect 1478 43488 1534 43544
rect 1602 43488 1658 43544
rect 1726 43488 1782 43544
rect 1850 43488 1906 43544
rect 114 43364 170 43420
rect 238 43364 294 43420
rect 362 43364 418 43420
rect 486 43364 542 43420
rect 610 43364 666 43420
rect 734 43364 790 43420
rect 858 43364 914 43420
rect 982 43364 1038 43420
rect 1106 43364 1162 43420
rect 1230 43364 1286 43420
rect 1354 43364 1410 43420
rect 1478 43364 1534 43420
rect 1602 43364 1658 43420
rect 1726 43364 1782 43420
rect 1850 43364 1906 43420
rect 114 43240 170 43296
rect 238 43240 294 43296
rect 362 43240 418 43296
rect 486 43240 542 43296
rect 610 43240 666 43296
rect 734 43240 790 43296
rect 858 43240 914 43296
rect 982 43240 1038 43296
rect 1106 43240 1162 43296
rect 1230 43240 1286 43296
rect 1354 43240 1410 43296
rect 1478 43240 1534 43296
rect 1602 43240 1658 43296
rect 1726 43240 1782 43296
rect 1850 43240 1906 43296
rect 114 43116 170 43172
rect 238 43116 294 43172
rect 362 43116 418 43172
rect 486 43116 542 43172
rect 610 43116 666 43172
rect 734 43116 790 43172
rect 858 43116 914 43172
rect 982 43116 1038 43172
rect 1106 43116 1162 43172
rect 1230 43116 1286 43172
rect 1354 43116 1410 43172
rect 1478 43116 1534 43172
rect 1602 43116 1658 43172
rect 1726 43116 1782 43172
rect 1850 43116 1906 43172
rect 114 42992 170 43048
rect 238 42992 294 43048
rect 362 42992 418 43048
rect 486 42992 542 43048
rect 610 42992 666 43048
rect 734 42992 790 43048
rect 858 42992 914 43048
rect 982 42992 1038 43048
rect 1106 42992 1162 43048
rect 1230 42992 1286 43048
rect 1354 42992 1410 43048
rect 1478 42992 1534 43048
rect 1602 42992 1658 43048
rect 1726 42992 1782 43048
rect 1850 42992 1906 43048
rect 114 42431 170 42487
rect 238 42431 294 42487
rect 362 42431 418 42487
rect 486 42431 542 42487
rect 610 42431 666 42487
rect 734 42431 790 42487
rect 858 42431 914 42487
rect 982 42431 1038 42487
rect 1106 42431 1162 42487
rect 1230 42431 1286 42487
rect 1354 42431 1410 42487
rect 1478 42431 1534 42487
rect 1602 42431 1658 42487
rect 1726 42431 1782 42487
rect 1850 42431 1906 42487
rect 114 42307 170 42363
rect 238 42307 294 42363
rect 362 42307 418 42363
rect 486 42307 542 42363
rect 610 42307 666 42363
rect 734 42307 790 42363
rect 858 42307 914 42363
rect 982 42307 1038 42363
rect 1106 42307 1162 42363
rect 1230 42307 1286 42363
rect 1354 42307 1410 42363
rect 1478 42307 1534 42363
rect 1602 42307 1658 42363
rect 1726 42307 1782 42363
rect 1850 42307 1906 42363
rect 114 42183 170 42239
rect 238 42183 294 42239
rect 362 42183 418 42239
rect 486 42183 542 42239
rect 610 42183 666 42239
rect 734 42183 790 42239
rect 858 42183 914 42239
rect 982 42183 1038 42239
rect 1106 42183 1162 42239
rect 1230 42183 1286 42239
rect 1354 42183 1410 42239
rect 1478 42183 1534 42239
rect 1602 42183 1658 42239
rect 1726 42183 1782 42239
rect 1850 42183 1906 42239
rect 114 42059 170 42115
rect 238 42059 294 42115
rect 362 42059 418 42115
rect 486 42059 542 42115
rect 610 42059 666 42115
rect 734 42059 790 42115
rect 858 42059 914 42115
rect 982 42059 1038 42115
rect 1106 42059 1162 42115
rect 1230 42059 1286 42115
rect 1354 42059 1410 42115
rect 1478 42059 1534 42115
rect 1602 42059 1658 42115
rect 1726 42059 1782 42115
rect 1850 42059 1906 42115
rect 114 41935 170 41991
rect 238 41935 294 41991
rect 362 41935 418 41991
rect 486 41935 542 41991
rect 610 41935 666 41991
rect 734 41935 790 41991
rect 858 41935 914 41991
rect 982 41935 1038 41991
rect 1106 41935 1162 41991
rect 1230 41935 1286 41991
rect 1354 41935 1410 41991
rect 1478 41935 1534 41991
rect 1602 41935 1658 41991
rect 1726 41935 1782 41991
rect 1850 41935 1906 41991
rect 114 41811 170 41867
rect 238 41811 294 41867
rect 362 41811 418 41867
rect 486 41811 542 41867
rect 610 41811 666 41867
rect 734 41811 790 41867
rect 858 41811 914 41867
rect 982 41811 1038 41867
rect 1106 41811 1162 41867
rect 1230 41811 1286 41867
rect 1354 41811 1410 41867
rect 1478 41811 1534 41867
rect 1602 41811 1658 41867
rect 1726 41811 1782 41867
rect 1850 41811 1906 41867
rect 114 41687 170 41743
rect 238 41687 294 41743
rect 362 41687 418 41743
rect 486 41687 542 41743
rect 610 41687 666 41743
rect 734 41687 790 41743
rect 858 41687 914 41743
rect 982 41687 1038 41743
rect 1106 41687 1162 41743
rect 1230 41687 1286 41743
rect 1354 41687 1410 41743
rect 1478 41687 1534 41743
rect 1602 41687 1658 41743
rect 1726 41687 1782 41743
rect 1850 41687 1906 41743
rect 114 41563 170 41619
rect 238 41563 294 41619
rect 362 41563 418 41619
rect 486 41563 542 41619
rect 610 41563 666 41619
rect 734 41563 790 41619
rect 858 41563 914 41619
rect 982 41563 1038 41619
rect 1106 41563 1162 41619
rect 1230 41563 1286 41619
rect 1354 41563 1410 41619
rect 1478 41563 1534 41619
rect 1602 41563 1658 41619
rect 1726 41563 1782 41619
rect 1850 41563 1906 41619
rect 114 41439 170 41495
rect 238 41439 294 41495
rect 362 41439 418 41495
rect 486 41439 542 41495
rect 610 41439 666 41495
rect 734 41439 790 41495
rect 858 41439 914 41495
rect 982 41439 1038 41495
rect 1106 41439 1162 41495
rect 1230 41439 1286 41495
rect 1354 41439 1410 41495
rect 1478 41439 1534 41495
rect 1602 41439 1658 41495
rect 1726 41439 1782 41495
rect 1850 41439 1906 41495
rect 114 41315 170 41371
rect 238 41315 294 41371
rect 362 41315 418 41371
rect 486 41315 542 41371
rect 610 41315 666 41371
rect 734 41315 790 41371
rect 858 41315 914 41371
rect 982 41315 1038 41371
rect 1106 41315 1162 41371
rect 1230 41315 1286 41371
rect 1354 41315 1410 41371
rect 1478 41315 1534 41371
rect 1602 41315 1658 41371
rect 1726 41315 1782 41371
rect 1850 41315 1906 41371
rect 114 40835 170 40891
rect 238 40835 294 40891
rect 362 40835 418 40891
rect 486 40835 542 40891
rect 610 40835 666 40891
rect 734 40835 790 40891
rect 858 40835 914 40891
rect 982 40835 1038 40891
rect 1106 40835 1162 40891
rect 1230 40835 1286 40891
rect 1354 40835 1410 40891
rect 1478 40835 1534 40891
rect 1602 40835 1658 40891
rect 1726 40835 1782 40891
rect 1850 40835 1906 40891
rect 114 40711 170 40767
rect 238 40711 294 40767
rect 362 40711 418 40767
rect 486 40711 542 40767
rect 610 40711 666 40767
rect 734 40711 790 40767
rect 858 40711 914 40767
rect 982 40711 1038 40767
rect 1106 40711 1162 40767
rect 1230 40711 1286 40767
rect 1354 40711 1410 40767
rect 1478 40711 1534 40767
rect 1602 40711 1658 40767
rect 1726 40711 1782 40767
rect 1850 40711 1906 40767
rect 114 40587 170 40643
rect 238 40587 294 40643
rect 362 40587 418 40643
rect 486 40587 542 40643
rect 610 40587 666 40643
rect 734 40587 790 40643
rect 858 40587 914 40643
rect 982 40587 1038 40643
rect 1106 40587 1162 40643
rect 1230 40587 1286 40643
rect 1354 40587 1410 40643
rect 1478 40587 1534 40643
rect 1602 40587 1658 40643
rect 1726 40587 1782 40643
rect 1850 40587 1906 40643
rect 114 40463 170 40519
rect 238 40463 294 40519
rect 362 40463 418 40519
rect 486 40463 542 40519
rect 610 40463 666 40519
rect 734 40463 790 40519
rect 858 40463 914 40519
rect 982 40463 1038 40519
rect 1106 40463 1162 40519
rect 1230 40463 1286 40519
rect 1354 40463 1410 40519
rect 1478 40463 1534 40519
rect 1602 40463 1658 40519
rect 1726 40463 1782 40519
rect 1850 40463 1906 40519
rect 114 40339 170 40395
rect 238 40339 294 40395
rect 362 40339 418 40395
rect 486 40339 542 40395
rect 610 40339 666 40395
rect 734 40339 790 40395
rect 858 40339 914 40395
rect 982 40339 1038 40395
rect 1106 40339 1162 40395
rect 1230 40339 1286 40395
rect 1354 40339 1410 40395
rect 1478 40339 1534 40395
rect 1602 40339 1658 40395
rect 1726 40339 1782 40395
rect 1850 40339 1906 40395
rect 114 40215 170 40271
rect 238 40215 294 40271
rect 362 40215 418 40271
rect 486 40215 542 40271
rect 610 40215 666 40271
rect 734 40215 790 40271
rect 858 40215 914 40271
rect 982 40215 1038 40271
rect 1106 40215 1162 40271
rect 1230 40215 1286 40271
rect 1354 40215 1410 40271
rect 1478 40215 1534 40271
rect 1602 40215 1658 40271
rect 1726 40215 1782 40271
rect 1850 40215 1906 40271
rect 114 40091 170 40147
rect 238 40091 294 40147
rect 362 40091 418 40147
rect 486 40091 542 40147
rect 610 40091 666 40147
rect 734 40091 790 40147
rect 858 40091 914 40147
rect 982 40091 1038 40147
rect 1106 40091 1162 40147
rect 1230 40091 1286 40147
rect 1354 40091 1410 40147
rect 1478 40091 1534 40147
rect 1602 40091 1658 40147
rect 1726 40091 1782 40147
rect 1850 40091 1906 40147
rect 114 39967 170 40023
rect 238 39967 294 40023
rect 362 39967 418 40023
rect 486 39967 542 40023
rect 610 39967 666 40023
rect 734 39967 790 40023
rect 858 39967 914 40023
rect 982 39967 1038 40023
rect 1106 39967 1162 40023
rect 1230 39967 1286 40023
rect 1354 39967 1410 40023
rect 1478 39967 1534 40023
rect 1602 39967 1658 40023
rect 1726 39967 1782 40023
rect 1850 39967 1906 40023
rect 114 39843 170 39899
rect 238 39843 294 39899
rect 362 39843 418 39899
rect 486 39843 542 39899
rect 610 39843 666 39899
rect 734 39843 790 39899
rect 858 39843 914 39899
rect 982 39843 1038 39899
rect 1106 39843 1162 39899
rect 1230 39843 1286 39899
rect 1354 39843 1410 39899
rect 1478 39843 1534 39899
rect 1602 39843 1658 39899
rect 1726 39843 1782 39899
rect 1850 39843 1906 39899
rect 114 39719 170 39775
rect 238 39719 294 39775
rect 362 39719 418 39775
rect 486 39719 542 39775
rect 610 39719 666 39775
rect 734 39719 790 39775
rect 858 39719 914 39775
rect 982 39719 1038 39775
rect 1106 39719 1162 39775
rect 1230 39719 1286 39775
rect 1354 39719 1410 39775
rect 1478 39719 1534 39775
rect 1602 39719 1658 39775
rect 1726 39719 1782 39775
rect 1850 39719 1906 39775
rect 114 39188 170 39244
rect 238 39188 294 39244
rect 362 39188 418 39244
rect 486 39188 542 39244
rect 610 39188 666 39244
rect 734 39188 790 39244
rect 858 39188 914 39244
rect 982 39188 1038 39244
rect 1106 39188 1162 39244
rect 1230 39188 1286 39244
rect 1354 39188 1410 39244
rect 1478 39188 1534 39244
rect 1602 39188 1658 39244
rect 1726 39188 1782 39244
rect 1850 39188 1906 39244
rect 114 39064 170 39120
rect 238 39064 294 39120
rect 362 39064 418 39120
rect 486 39064 542 39120
rect 610 39064 666 39120
rect 734 39064 790 39120
rect 858 39064 914 39120
rect 982 39064 1038 39120
rect 1106 39064 1162 39120
rect 1230 39064 1286 39120
rect 1354 39064 1410 39120
rect 1478 39064 1534 39120
rect 1602 39064 1658 39120
rect 1726 39064 1782 39120
rect 1850 39064 1906 39120
rect 114 38940 170 38996
rect 238 38940 294 38996
rect 362 38940 418 38996
rect 486 38940 542 38996
rect 610 38940 666 38996
rect 734 38940 790 38996
rect 858 38940 914 38996
rect 982 38940 1038 38996
rect 1106 38940 1162 38996
rect 1230 38940 1286 38996
rect 1354 38940 1410 38996
rect 1478 38940 1534 38996
rect 1602 38940 1658 38996
rect 1726 38940 1782 38996
rect 1850 38940 1906 38996
rect 114 38816 170 38872
rect 238 38816 294 38872
rect 362 38816 418 38872
rect 486 38816 542 38872
rect 610 38816 666 38872
rect 734 38816 790 38872
rect 858 38816 914 38872
rect 982 38816 1038 38872
rect 1106 38816 1162 38872
rect 1230 38816 1286 38872
rect 1354 38816 1410 38872
rect 1478 38816 1534 38872
rect 1602 38816 1658 38872
rect 1726 38816 1782 38872
rect 1850 38816 1906 38872
rect 114 38692 170 38748
rect 238 38692 294 38748
rect 362 38692 418 38748
rect 486 38692 542 38748
rect 610 38692 666 38748
rect 734 38692 790 38748
rect 858 38692 914 38748
rect 982 38692 1038 38748
rect 1106 38692 1162 38748
rect 1230 38692 1286 38748
rect 1354 38692 1410 38748
rect 1478 38692 1534 38748
rect 1602 38692 1658 38748
rect 1726 38692 1782 38748
rect 1850 38692 1906 38748
rect 114 38568 170 38624
rect 238 38568 294 38624
rect 362 38568 418 38624
rect 486 38568 542 38624
rect 610 38568 666 38624
rect 734 38568 790 38624
rect 858 38568 914 38624
rect 982 38568 1038 38624
rect 1106 38568 1162 38624
rect 1230 38568 1286 38624
rect 1354 38568 1410 38624
rect 1478 38568 1534 38624
rect 1602 38568 1658 38624
rect 1726 38568 1782 38624
rect 1850 38568 1906 38624
rect 114 38444 170 38500
rect 238 38444 294 38500
rect 362 38444 418 38500
rect 486 38444 542 38500
rect 610 38444 666 38500
rect 734 38444 790 38500
rect 858 38444 914 38500
rect 982 38444 1038 38500
rect 1106 38444 1162 38500
rect 1230 38444 1286 38500
rect 1354 38444 1410 38500
rect 1478 38444 1534 38500
rect 1602 38444 1658 38500
rect 1726 38444 1782 38500
rect 1850 38444 1906 38500
rect 114 38320 170 38376
rect 238 38320 294 38376
rect 362 38320 418 38376
rect 486 38320 542 38376
rect 610 38320 666 38376
rect 734 38320 790 38376
rect 858 38320 914 38376
rect 982 38320 1038 38376
rect 1106 38320 1162 38376
rect 1230 38320 1286 38376
rect 1354 38320 1410 38376
rect 1478 38320 1534 38376
rect 1602 38320 1658 38376
rect 1726 38320 1782 38376
rect 1850 38320 1906 38376
rect 114 38196 170 38252
rect 238 38196 294 38252
rect 362 38196 418 38252
rect 486 38196 542 38252
rect 610 38196 666 38252
rect 734 38196 790 38252
rect 858 38196 914 38252
rect 982 38196 1038 38252
rect 1106 38196 1162 38252
rect 1230 38196 1286 38252
rect 1354 38196 1410 38252
rect 1478 38196 1534 38252
rect 1602 38196 1658 38252
rect 1726 38196 1782 38252
rect 1850 38196 1906 38252
rect 114 38072 170 38128
rect 238 38072 294 38128
rect 362 38072 418 38128
rect 486 38072 542 38128
rect 610 38072 666 38128
rect 734 38072 790 38128
rect 858 38072 914 38128
rect 982 38072 1038 38128
rect 1106 38072 1162 38128
rect 1230 38072 1286 38128
rect 1354 38072 1410 38128
rect 1478 38072 1534 38128
rect 1602 38072 1658 38128
rect 1726 38072 1782 38128
rect 1850 38072 1906 38128
rect 114 37948 170 38004
rect 238 37948 294 38004
rect 362 37948 418 38004
rect 486 37948 542 38004
rect 610 37948 666 38004
rect 734 37948 790 38004
rect 858 37948 914 38004
rect 982 37948 1038 38004
rect 1106 37948 1162 38004
rect 1230 37948 1286 38004
rect 1354 37948 1410 38004
rect 1478 37948 1534 38004
rect 1602 37948 1658 38004
rect 1726 37948 1782 38004
rect 1850 37948 1906 38004
rect 114 37824 170 37880
rect 238 37824 294 37880
rect 362 37824 418 37880
rect 486 37824 542 37880
rect 610 37824 666 37880
rect 734 37824 790 37880
rect 858 37824 914 37880
rect 982 37824 1038 37880
rect 1106 37824 1162 37880
rect 1230 37824 1286 37880
rect 1354 37824 1410 37880
rect 1478 37824 1534 37880
rect 1602 37824 1658 37880
rect 1726 37824 1782 37880
rect 1850 37824 1906 37880
rect 114 37700 170 37756
rect 238 37700 294 37756
rect 362 37700 418 37756
rect 486 37700 542 37756
rect 610 37700 666 37756
rect 734 37700 790 37756
rect 858 37700 914 37756
rect 982 37700 1038 37756
rect 1106 37700 1162 37756
rect 1230 37700 1286 37756
rect 1354 37700 1410 37756
rect 1478 37700 1534 37756
rect 1602 37700 1658 37756
rect 1726 37700 1782 37756
rect 1850 37700 1906 37756
rect 114 37576 170 37632
rect 238 37576 294 37632
rect 362 37576 418 37632
rect 486 37576 542 37632
rect 610 37576 666 37632
rect 734 37576 790 37632
rect 858 37576 914 37632
rect 982 37576 1038 37632
rect 1106 37576 1162 37632
rect 1230 37576 1286 37632
rect 1354 37576 1410 37632
rect 1478 37576 1534 37632
rect 1602 37576 1658 37632
rect 1726 37576 1782 37632
rect 1850 37576 1906 37632
rect 114 37452 170 37508
rect 238 37452 294 37508
rect 362 37452 418 37508
rect 486 37452 542 37508
rect 610 37452 666 37508
rect 734 37452 790 37508
rect 858 37452 914 37508
rect 982 37452 1038 37508
rect 1106 37452 1162 37508
rect 1230 37452 1286 37508
rect 1354 37452 1410 37508
rect 1478 37452 1534 37508
rect 1602 37452 1658 37508
rect 1726 37452 1782 37508
rect 1850 37452 1906 37508
rect 114 37328 170 37384
rect 238 37328 294 37384
rect 362 37328 418 37384
rect 486 37328 542 37384
rect 610 37328 666 37384
rect 734 37328 790 37384
rect 858 37328 914 37384
rect 982 37328 1038 37384
rect 1106 37328 1162 37384
rect 1230 37328 1286 37384
rect 1354 37328 1410 37384
rect 1478 37328 1534 37384
rect 1602 37328 1658 37384
rect 1726 37328 1782 37384
rect 1850 37328 1906 37384
rect 114 37204 170 37260
rect 238 37204 294 37260
rect 362 37204 418 37260
rect 486 37204 542 37260
rect 610 37204 666 37260
rect 734 37204 790 37260
rect 858 37204 914 37260
rect 982 37204 1038 37260
rect 1106 37204 1162 37260
rect 1230 37204 1286 37260
rect 1354 37204 1410 37260
rect 1478 37204 1534 37260
rect 1602 37204 1658 37260
rect 1726 37204 1782 37260
rect 1850 37204 1906 37260
rect 114 37080 170 37136
rect 238 37080 294 37136
rect 362 37080 418 37136
rect 486 37080 542 37136
rect 610 37080 666 37136
rect 734 37080 790 37136
rect 858 37080 914 37136
rect 982 37080 1038 37136
rect 1106 37080 1162 37136
rect 1230 37080 1286 37136
rect 1354 37080 1410 37136
rect 1478 37080 1534 37136
rect 1602 37080 1658 37136
rect 1726 37080 1782 37136
rect 1850 37080 1906 37136
rect 114 36956 170 37012
rect 238 36956 294 37012
rect 362 36956 418 37012
rect 486 36956 542 37012
rect 610 36956 666 37012
rect 734 36956 790 37012
rect 858 36956 914 37012
rect 982 36956 1038 37012
rect 1106 36956 1162 37012
rect 1230 36956 1286 37012
rect 1354 36956 1410 37012
rect 1478 36956 1534 37012
rect 1602 36956 1658 37012
rect 1726 36956 1782 37012
rect 1850 36956 1906 37012
rect 114 36832 170 36888
rect 238 36832 294 36888
rect 362 36832 418 36888
rect 486 36832 542 36888
rect 610 36832 666 36888
rect 734 36832 790 36888
rect 858 36832 914 36888
rect 982 36832 1038 36888
rect 1106 36832 1162 36888
rect 1230 36832 1286 36888
rect 1354 36832 1410 36888
rect 1478 36832 1534 36888
rect 1602 36832 1658 36888
rect 1726 36832 1782 36888
rect 1850 36832 1906 36888
rect 114 36708 170 36764
rect 238 36708 294 36764
rect 362 36708 418 36764
rect 486 36708 542 36764
rect 610 36708 666 36764
rect 734 36708 790 36764
rect 858 36708 914 36764
rect 982 36708 1038 36764
rect 1106 36708 1162 36764
rect 1230 36708 1286 36764
rect 1354 36708 1410 36764
rect 1478 36708 1534 36764
rect 1602 36708 1658 36764
rect 1726 36708 1782 36764
rect 1850 36708 1906 36764
rect 114 36584 170 36640
rect 238 36584 294 36640
rect 362 36584 418 36640
rect 486 36584 542 36640
rect 610 36584 666 36640
rect 734 36584 790 36640
rect 858 36584 914 36640
rect 982 36584 1038 36640
rect 1106 36584 1162 36640
rect 1230 36584 1286 36640
rect 1354 36584 1410 36640
rect 1478 36584 1534 36640
rect 1602 36584 1658 36640
rect 1726 36584 1782 36640
rect 1850 36584 1906 36640
rect 114 36003 170 36059
rect 238 36003 294 36059
rect 362 36003 418 36059
rect 486 36003 542 36059
rect 610 36003 666 36059
rect 734 36003 790 36059
rect 858 36003 914 36059
rect 982 36003 1038 36059
rect 1106 36003 1162 36059
rect 1230 36003 1286 36059
rect 1354 36003 1410 36059
rect 1478 36003 1534 36059
rect 1602 36003 1658 36059
rect 1726 36003 1782 36059
rect 1850 36003 1906 36059
rect 114 35879 170 35935
rect 238 35879 294 35935
rect 362 35879 418 35935
rect 486 35879 542 35935
rect 610 35879 666 35935
rect 734 35879 790 35935
rect 858 35879 914 35935
rect 982 35879 1038 35935
rect 1106 35879 1162 35935
rect 1230 35879 1286 35935
rect 1354 35879 1410 35935
rect 1478 35879 1534 35935
rect 1602 35879 1658 35935
rect 1726 35879 1782 35935
rect 1850 35879 1906 35935
rect 114 35755 170 35811
rect 238 35755 294 35811
rect 362 35755 418 35811
rect 486 35755 542 35811
rect 610 35755 666 35811
rect 734 35755 790 35811
rect 858 35755 914 35811
rect 982 35755 1038 35811
rect 1106 35755 1162 35811
rect 1230 35755 1286 35811
rect 1354 35755 1410 35811
rect 1478 35755 1534 35811
rect 1602 35755 1658 35811
rect 1726 35755 1782 35811
rect 1850 35755 1906 35811
rect 114 35631 170 35687
rect 238 35631 294 35687
rect 362 35631 418 35687
rect 486 35631 542 35687
rect 610 35631 666 35687
rect 734 35631 790 35687
rect 858 35631 914 35687
rect 982 35631 1038 35687
rect 1106 35631 1162 35687
rect 1230 35631 1286 35687
rect 1354 35631 1410 35687
rect 1478 35631 1534 35687
rect 1602 35631 1658 35687
rect 1726 35631 1782 35687
rect 1850 35631 1906 35687
rect 114 35507 170 35563
rect 238 35507 294 35563
rect 362 35507 418 35563
rect 486 35507 542 35563
rect 610 35507 666 35563
rect 734 35507 790 35563
rect 858 35507 914 35563
rect 982 35507 1038 35563
rect 1106 35507 1162 35563
rect 1230 35507 1286 35563
rect 1354 35507 1410 35563
rect 1478 35507 1534 35563
rect 1602 35507 1658 35563
rect 1726 35507 1782 35563
rect 1850 35507 1906 35563
rect 114 35383 170 35439
rect 238 35383 294 35439
rect 362 35383 418 35439
rect 486 35383 542 35439
rect 610 35383 666 35439
rect 734 35383 790 35439
rect 858 35383 914 35439
rect 982 35383 1038 35439
rect 1106 35383 1162 35439
rect 1230 35383 1286 35439
rect 1354 35383 1410 35439
rect 1478 35383 1534 35439
rect 1602 35383 1658 35439
rect 1726 35383 1782 35439
rect 1850 35383 1906 35439
rect 114 35259 170 35315
rect 238 35259 294 35315
rect 362 35259 418 35315
rect 486 35259 542 35315
rect 610 35259 666 35315
rect 734 35259 790 35315
rect 858 35259 914 35315
rect 982 35259 1038 35315
rect 1106 35259 1162 35315
rect 1230 35259 1286 35315
rect 1354 35259 1410 35315
rect 1478 35259 1534 35315
rect 1602 35259 1658 35315
rect 1726 35259 1782 35315
rect 1850 35259 1906 35315
rect 114 35135 170 35191
rect 238 35135 294 35191
rect 362 35135 418 35191
rect 486 35135 542 35191
rect 610 35135 666 35191
rect 734 35135 790 35191
rect 858 35135 914 35191
rect 982 35135 1038 35191
rect 1106 35135 1162 35191
rect 1230 35135 1286 35191
rect 1354 35135 1410 35191
rect 1478 35135 1534 35191
rect 1602 35135 1658 35191
rect 1726 35135 1782 35191
rect 1850 35135 1906 35191
rect 114 35011 170 35067
rect 238 35011 294 35067
rect 362 35011 418 35067
rect 486 35011 542 35067
rect 610 35011 666 35067
rect 734 35011 790 35067
rect 858 35011 914 35067
rect 982 35011 1038 35067
rect 1106 35011 1162 35067
rect 1230 35011 1286 35067
rect 1354 35011 1410 35067
rect 1478 35011 1534 35067
rect 1602 35011 1658 35067
rect 1726 35011 1782 35067
rect 1850 35011 1906 35067
rect 114 34887 170 34943
rect 238 34887 294 34943
rect 362 34887 418 34943
rect 486 34887 542 34943
rect 610 34887 666 34943
rect 734 34887 790 34943
rect 858 34887 914 34943
rect 982 34887 1038 34943
rect 1106 34887 1162 34943
rect 1230 34887 1286 34943
rect 1354 34887 1410 34943
rect 1478 34887 1534 34943
rect 1602 34887 1658 34943
rect 1726 34887 1782 34943
rect 1850 34887 1906 34943
rect 114 34763 170 34819
rect 238 34763 294 34819
rect 362 34763 418 34819
rect 486 34763 542 34819
rect 610 34763 666 34819
rect 734 34763 790 34819
rect 858 34763 914 34819
rect 982 34763 1038 34819
rect 1106 34763 1162 34819
rect 1230 34763 1286 34819
rect 1354 34763 1410 34819
rect 1478 34763 1534 34819
rect 1602 34763 1658 34819
rect 1726 34763 1782 34819
rect 1850 34763 1906 34819
rect 114 34639 170 34695
rect 238 34639 294 34695
rect 362 34639 418 34695
rect 486 34639 542 34695
rect 610 34639 666 34695
rect 734 34639 790 34695
rect 858 34639 914 34695
rect 982 34639 1038 34695
rect 1106 34639 1162 34695
rect 1230 34639 1286 34695
rect 1354 34639 1410 34695
rect 1478 34639 1534 34695
rect 1602 34639 1658 34695
rect 1726 34639 1782 34695
rect 1850 34639 1906 34695
rect 114 34515 170 34571
rect 238 34515 294 34571
rect 362 34515 418 34571
rect 486 34515 542 34571
rect 610 34515 666 34571
rect 734 34515 790 34571
rect 858 34515 914 34571
rect 982 34515 1038 34571
rect 1106 34515 1162 34571
rect 1230 34515 1286 34571
rect 1354 34515 1410 34571
rect 1478 34515 1534 34571
rect 1602 34515 1658 34571
rect 1726 34515 1782 34571
rect 1850 34515 1906 34571
rect 114 34391 170 34447
rect 238 34391 294 34447
rect 362 34391 418 34447
rect 486 34391 542 34447
rect 610 34391 666 34447
rect 734 34391 790 34447
rect 858 34391 914 34447
rect 982 34391 1038 34447
rect 1106 34391 1162 34447
rect 1230 34391 1286 34447
rect 1354 34391 1410 34447
rect 1478 34391 1534 34447
rect 1602 34391 1658 34447
rect 1726 34391 1782 34447
rect 1850 34391 1906 34447
rect 114 34267 170 34323
rect 238 34267 294 34323
rect 362 34267 418 34323
rect 486 34267 542 34323
rect 610 34267 666 34323
rect 734 34267 790 34323
rect 858 34267 914 34323
rect 982 34267 1038 34323
rect 1106 34267 1162 34323
rect 1230 34267 1286 34323
rect 1354 34267 1410 34323
rect 1478 34267 1534 34323
rect 1602 34267 1658 34323
rect 1726 34267 1782 34323
rect 1850 34267 1906 34323
rect 114 34143 170 34199
rect 238 34143 294 34199
rect 362 34143 418 34199
rect 486 34143 542 34199
rect 610 34143 666 34199
rect 734 34143 790 34199
rect 858 34143 914 34199
rect 982 34143 1038 34199
rect 1106 34143 1162 34199
rect 1230 34143 1286 34199
rect 1354 34143 1410 34199
rect 1478 34143 1534 34199
rect 1602 34143 1658 34199
rect 1726 34143 1782 34199
rect 1850 34143 1906 34199
rect 114 34019 170 34075
rect 238 34019 294 34075
rect 362 34019 418 34075
rect 486 34019 542 34075
rect 610 34019 666 34075
rect 734 34019 790 34075
rect 858 34019 914 34075
rect 982 34019 1038 34075
rect 1106 34019 1162 34075
rect 1230 34019 1286 34075
rect 1354 34019 1410 34075
rect 1478 34019 1534 34075
rect 1602 34019 1658 34075
rect 1726 34019 1782 34075
rect 1850 34019 1906 34075
rect 114 33895 170 33951
rect 238 33895 294 33951
rect 362 33895 418 33951
rect 486 33895 542 33951
rect 610 33895 666 33951
rect 734 33895 790 33951
rect 858 33895 914 33951
rect 982 33895 1038 33951
rect 1106 33895 1162 33951
rect 1230 33895 1286 33951
rect 1354 33895 1410 33951
rect 1478 33895 1534 33951
rect 1602 33895 1658 33951
rect 1726 33895 1782 33951
rect 1850 33895 1906 33951
rect 114 33771 170 33827
rect 238 33771 294 33827
rect 362 33771 418 33827
rect 486 33771 542 33827
rect 610 33771 666 33827
rect 734 33771 790 33827
rect 858 33771 914 33827
rect 982 33771 1038 33827
rect 1106 33771 1162 33827
rect 1230 33771 1286 33827
rect 1354 33771 1410 33827
rect 1478 33771 1534 33827
rect 1602 33771 1658 33827
rect 1726 33771 1782 33827
rect 1850 33771 1906 33827
rect 114 33647 170 33703
rect 238 33647 294 33703
rect 362 33647 418 33703
rect 486 33647 542 33703
rect 610 33647 666 33703
rect 734 33647 790 33703
rect 858 33647 914 33703
rect 982 33647 1038 33703
rect 1106 33647 1162 33703
rect 1230 33647 1286 33703
rect 1354 33647 1410 33703
rect 1478 33647 1534 33703
rect 1602 33647 1658 33703
rect 1726 33647 1782 33703
rect 1850 33647 1906 33703
rect 114 33523 170 33579
rect 238 33523 294 33579
rect 362 33523 418 33579
rect 486 33523 542 33579
rect 610 33523 666 33579
rect 734 33523 790 33579
rect 858 33523 914 33579
rect 982 33523 1038 33579
rect 1106 33523 1162 33579
rect 1230 33523 1286 33579
rect 1354 33523 1410 33579
rect 1478 33523 1534 33579
rect 1602 33523 1658 33579
rect 1726 33523 1782 33579
rect 1850 33523 1906 33579
rect 114 33399 170 33455
rect 238 33399 294 33455
rect 362 33399 418 33455
rect 486 33399 542 33455
rect 610 33399 666 33455
rect 734 33399 790 33455
rect 858 33399 914 33455
rect 982 33399 1038 33455
rect 1106 33399 1162 33455
rect 1230 33399 1286 33455
rect 1354 33399 1410 33455
rect 1478 33399 1534 33455
rect 1602 33399 1658 33455
rect 1726 33399 1782 33455
rect 1850 33399 1906 33455
rect 114 32788 170 32844
rect 238 32788 294 32844
rect 362 32788 418 32844
rect 486 32788 542 32844
rect 610 32788 666 32844
rect 734 32788 790 32844
rect 858 32788 914 32844
rect 982 32788 1038 32844
rect 1106 32788 1162 32844
rect 1230 32788 1286 32844
rect 1354 32788 1410 32844
rect 1478 32788 1534 32844
rect 1602 32788 1658 32844
rect 1726 32788 1782 32844
rect 1850 32788 1906 32844
rect 114 32664 170 32720
rect 238 32664 294 32720
rect 362 32664 418 32720
rect 486 32664 542 32720
rect 610 32664 666 32720
rect 734 32664 790 32720
rect 858 32664 914 32720
rect 982 32664 1038 32720
rect 1106 32664 1162 32720
rect 1230 32664 1286 32720
rect 1354 32664 1410 32720
rect 1478 32664 1534 32720
rect 1602 32664 1658 32720
rect 1726 32664 1782 32720
rect 1850 32664 1906 32720
rect 114 32540 170 32596
rect 238 32540 294 32596
rect 362 32540 418 32596
rect 486 32540 542 32596
rect 610 32540 666 32596
rect 734 32540 790 32596
rect 858 32540 914 32596
rect 982 32540 1038 32596
rect 1106 32540 1162 32596
rect 1230 32540 1286 32596
rect 1354 32540 1410 32596
rect 1478 32540 1534 32596
rect 1602 32540 1658 32596
rect 1726 32540 1782 32596
rect 1850 32540 1906 32596
rect 114 32416 170 32472
rect 238 32416 294 32472
rect 362 32416 418 32472
rect 486 32416 542 32472
rect 610 32416 666 32472
rect 734 32416 790 32472
rect 858 32416 914 32472
rect 982 32416 1038 32472
rect 1106 32416 1162 32472
rect 1230 32416 1286 32472
rect 1354 32416 1410 32472
rect 1478 32416 1534 32472
rect 1602 32416 1658 32472
rect 1726 32416 1782 32472
rect 1850 32416 1906 32472
rect 114 32292 170 32348
rect 238 32292 294 32348
rect 362 32292 418 32348
rect 486 32292 542 32348
rect 610 32292 666 32348
rect 734 32292 790 32348
rect 858 32292 914 32348
rect 982 32292 1038 32348
rect 1106 32292 1162 32348
rect 1230 32292 1286 32348
rect 1354 32292 1410 32348
rect 1478 32292 1534 32348
rect 1602 32292 1658 32348
rect 1726 32292 1782 32348
rect 1850 32292 1906 32348
rect 114 32168 170 32224
rect 238 32168 294 32224
rect 362 32168 418 32224
rect 486 32168 542 32224
rect 610 32168 666 32224
rect 734 32168 790 32224
rect 858 32168 914 32224
rect 982 32168 1038 32224
rect 1106 32168 1162 32224
rect 1230 32168 1286 32224
rect 1354 32168 1410 32224
rect 1478 32168 1534 32224
rect 1602 32168 1658 32224
rect 1726 32168 1782 32224
rect 1850 32168 1906 32224
rect 114 32044 170 32100
rect 238 32044 294 32100
rect 362 32044 418 32100
rect 486 32044 542 32100
rect 610 32044 666 32100
rect 734 32044 790 32100
rect 858 32044 914 32100
rect 982 32044 1038 32100
rect 1106 32044 1162 32100
rect 1230 32044 1286 32100
rect 1354 32044 1410 32100
rect 1478 32044 1534 32100
rect 1602 32044 1658 32100
rect 1726 32044 1782 32100
rect 1850 32044 1906 32100
rect 114 31920 170 31976
rect 238 31920 294 31976
rect 362 31920 418 31976
rect 486 31920 542 31976
rect 610 31920 666 31976
rect 734 31920 790 31976
rect 858 31920 914 31976
rect 982 31920 1038 31976
rect 1106 31920 1162 31976
rect 1230 31920 1286 31976
rect 1354 31920 1410 31976
rect 1478 31920 1534 31976
rect 1602 31920 1658 31976
rect 1726 31920 1782 31976
rect 1850 31920 1906 31976
rect 114 31796 170 31852
rect 238 31796 294 31852
rect 362 31796 418 31852
rect 486 31796 542 31852
rect 610 31796 666 31852
rect 734 31796 790 31852
rect 858 31796 914 31852
rect 982 31796 1038 31852
rect 1106 31796 1162 31852
rect 1230 31796 1286 31852
rect 1354 31796 1410 31852
rect 1478 31796 1534 31852
rect 1602 31796 1658 31852
rect 1726 31796 1782 31852
rect 1850 31796 1906 31852
rect 114 31672 170 31728
rect 238 31672 294 31728
rect 362 31672 418 31728
rect 486 31672 542 31728
rect 610 31672 666 31728
rect 734 31672 790 31728
rect 858 31672 914 31728
rect 982 31672 1038 31728
rect 1106 31672 1162 31728
rect 1230 31672 1286 31728
rect 1354 31672 1410 31728
rect 1478 31672 1534 31728
rect 1602 31672 1658 31728
rect 1726 31672 1782 31728
rect 1850 31672 1906 31728
rect 114 31548 170 31604
rect 238 31548 294 31604
rect 362 31548 418 31604
rect 486 31548 542 31604
rect 610 31548 666 31604
rect 734 31548 790 31604
rect 858 31548 914 31604
rect 982 31548 1038 31604
rect 1106 31548 1162 31604
rect 1230 31548 1286 31604
rect 1354 31548 1410 31604
rect 1478 31548 1534 31604
rect 1602 31548 1658 31604
rect 1726 31548 1782 31604
rect 1850 31548 1906 31604
rect 114 31424 170 31480
rect 238 31424 294 31480
rect 362 31424 418 31480
rect 486 31424 542 31480
rect 610 31424 666 31480
rect 734 31424 790 31480
rect 858 31424 914 31480
rect 982 31424 1038 31480
rect 1106 31424 1162 31480
rect 1230 31424 1286 31480
rect 1354 31424 1410 31480
rect 1478 31424 1534 31480
rect 1602 31424 1658 31480
rect 1726 31424 1782 31480
rect 1850 31424 1906 31480
rect 114 31300 170 31356
rect 238 31300 294 31356
rect 362 31300 418 31356
rect 486 31300 542 31356
rect 610 31300 666 31356
rect 734 31300 790 31356
rect 858 31300 914 31356
rect 982 31300 1038 31356
rect 1106 31300 1162 31356
rect 1230 31300 1286 31356
rect 1354 31300 1410 31356
rect 1478 31300 1534 31356
rect 1602 31300 1658 31356
rect 1726 31300 1782 31356
rect 1850 31300 1906 31356
rect 114 31176 170 31232
rect 238 31176 294 31232
rect 362 31176 418 31232
rect 486 31176 542 31232
rect 610 31176 666 31232
rect 734 31176 790 31232
rect 858 31176 914 31232
rect 982 31176 1038 31232
rect 1106 31176 1162 31232
rect 1230 31176 1286 31232
rect 1354 31176 1410 31232
rect 1478 31176 1534 31232
rect 1602 31176 1658 31232
rect 1726 31176 1782 31232
rect 1850 31176 1906 31232
rect 114 31052 170 31108
rect 238 31052 294 31108
rect 362 31052 418 31108
rect 486 31052 542 31108
rect 610 31052 666 31108
rect 734 31052 790 31108
rect 858 31052 914 31108
rect 982 31052 1038 31108
rect 1106 31052 1162 31108
rect 1230 31052 1286 31108
rect 1354 31052 1410 31108
rect 1478 31052 1534 31108
rect 1602 31052 1658 31108
rect 1726 31052 1782 31108
rect 1850 31052 1906 31108
rect 114 30928 170 30984
rect 238 30928 294 30984
rect 362 30928 418 30984
rect 486 30928 542 30984
rect 610 30928 666 30984
rect 734 30928 790 30984
rect 858 30928 914 30984
rect 982 30928 1038 30984
rect 1106 30928 1162 30984
rect 1230 30928 1286 30984
rect 1354 30928 1410 30984
rect 1478 30928 1534 30984
rect 1602 30928 1658 30984
rect 1726 30928 1782 30984
rect 1850 30928 1906 30984
rect 114 30804 170 30860
rect 238 30804 294 30860
rect 362 30804 418 30860
rect 486 30804 542 30860
rect 610 30804 666 30860
rect 734 30804 790 30860
rect 858 30804 914 30860
rect 982 30804 1038 30860
rect 1106 30804 1162 30860
rect 1230 30804 1286 30860
rect 1354 30804 1410 30860
rect 1478 30804 1534 30860
rect 1602 30804 1658 30860
rect 1726 30804 1782 30860
rect 1850 30804 1906 30860
rect 114 30680 170 30736
rect 238 30680 294 30736
rect 362 30680 418 30736
rect 486 30680 542 30736
rect 610 30680 666 30736
rect 734 30680 790 30736
rect 858 30680 914 30736
rect 982 30680 1038 30736
rect 1106 30680 1162 30736
rect 1230 30680 1286 30736
rect 1354 30680 1410 30736
rect 1478 30680 1534 30736
rect 1602 30680 1658 30736
rect 1726 30680 1782 30736
rect 1850 30680 1906 30736
rect 114 30556 170 30612
rect 238 30556 294 30612
rect 362 30556 418 30612
rect 486 30556 542 30612
rect 610 30556 666 30612
rect 734 30556 790 30612
rect 858 30556 914 30612
rect 982 30556 1038 30612
rect 1106 30556 1162 30612
rect 1230 30556 1286 30612
rect 1354 30556 1410 30612
rect 1478 30556 1534 30612
rect 1602 30556 1658 30612
rect 1726 30556 1782 30612
rect 1850 30556 1906 30612
rect 114 30432 170 30488
rect 238 30432 294 30488
rect 362 30432 418 30488
rect 486 30432 542 30488
rect 610 30432 666 30488
rect 734 30432 790 30488
rect 858 30432 914 30488
rect 982 30432 1038 30488
rect 1106 30432 1162 30488
rect 1230 30432 1286 30488
rect 1354 30432 1410 30488
rect 1478 30432 1534 30488
rect 1602 30432 1658 30488
rect 1726 30432 1782 30488
rect 1850 30432 1906 30488
rect 114 30308 170 30364
rect 238 30308 294 30364
rect 362 30308 418 30364
rect 486 30308 542 30364
rect 610 30308 666 30364
rect 734 30308 790 30364
rect 858 30308 914 30364
rect 982 30308 1038 30364
rect 1106 30308 1162 30364
rect 1230 30308 1286 30364
rect 1354 30308 1410 30364
rect 1478 30308 1534 30364
rect 1602 30308 1658 30364
rect 1726 30308 1782 30364
rect 1850 30308 1906 30364
rect 114 30184 170 30240
rect 238 30184 294 30240
rect 362 30184 418 30240
rect 486 30184 542 30240
rect 610 30184 666 30240
rect 734 30184 790 30240
rect 858 30184 914 30240
rect 982 30184 1038 30240
rect 1106 30184 1162 30240
rect 1230 30184 1286 30240
rect 1354 30184 1410 30240
rect 1478 30184 1534 30240
rect 1602 30184 1658 30240
rect 1726 30184 1782 30240
rect 1850 30184 1906 30240
rect 114 29587 170 29643
rect 238 29587 294 29643
rect 362 29587 418 29643
rect 486 29587 542 29643
rect 610 29587 666 29643
rect 734 29587 790 29643
rect 858 29587 914 29643
rect 982 29587 1038 29643
rect 1106 29587 1162 29643
rect 1230 29587 1286 29643
rect 1354 29587 1410 29643
rect 1478 29587 1534 29643
rect 1602 29587 1658 29643
rect 1726 29587 1782 29643
rect 1850 29587 1906 29643
rect 114 29463 170 29519
rect 238 29463 294 29519
rect 362 29463 418 29519
rect 486 29463 542 29519
rect 610 29463 666 29519
rect 734 29463 790 29519
rect 858 29463 914 29519
rect 982 29463 1038 29519
rect 1106 29463 1162 29519
rect 1230 29463 1286 29519
rect 1354 29463 1410 29519
rect 1478 29463 1534 29519
rect 1602 29463 1658 29519
rect 1726 29463 1782 29519
rect 1850 29463 1906 29519
rect 114 29339 170 29395
rect 238 29339 294 29395
rect 362 29339 418 29395
rect 486 29339 542 29395
rect 610 29339 666 29395
rect 734 29339 790 29395
rect 858 29339 914 29395
rect 982 29339 1038 29395
rect 1106 29339 1162 29395
rect 1230 29339 1286 29395
rect 1354 29339 1410 29395
rect 1478 29339 1534 29395
rect 1602 29339 1658 29395
rect 1726 29339 1782 29395
rect 1850 29339 1906 29395
rect 114 29215 170 29271
rect 238 29215 294 29271
rect 362 29215 418 29271
rect 486 29215 542 29271
rect 610 29215 666 29271
rect 734 29215 790 29271
rect 858 29215 914 29271
rect 982 29215 1038 29271
rect 1106 29215 1162 29271
rect 1230 29215 1286 29271
rect 1354 29215 1410 29271
rect 1478 29215 1534 29271
rect 1602 29215 1658 29271
rect 1726 29215 1782 29271
rect 1850 29215 1906 29271
rect 114 29091 170 29147
rect 238 29091 294 29147
rect 362 29091 418 29147
rect 486 29091 542 29147
rect 610 29091 666 29147
rect 734 29091 790 29147
rect 858 29091 914 29147
rect 982 29091 1038 29147
rect 1106 29091 1162 29147
rect 1230 29091 1286 29147
rect 1354 29091 1410 29147
rect 1478 29091 1534 29147
rect 1602 29091 1658 29147
rect 1726 29091 1782 29147
rect 1850 29091 1906 29147
rect 114 28967 170 29023
rect 238 28967 294 29023
rect 362 28967 418 29023
rect 486 28967 542 29023
rect 610 28967 666 29023
rect 734 28967 790 29023
rect 858 28967 914 29023
rect 982 28967 1038 29023
rect 1106 28967 1162 29023
rect 1230 28967 1286 29023
rect 1354 28967 1410 29023
rect 1478 28967 1534 29023
rect 1602 28967 1658 29023
rect 1726 28967 1782 29023
rect 1850 28967 1906 29023
rect 114 28843 170 28899
rect 238 28843 294 28899
rect 362 28843 418 28899
rect 486 28843 542 28899
rect 610 28843 666 28899
rect 734 28843 790 28899
rect 858 28843 914 28899
rect 982 28843 1038 28899
rect 1106 28843 1162 28899
rect 1230 28843 1286 28899
rect 1354 28843 1410 28899
rect 1478 28843 1534 28899
rect 1602 28843 1658 28899
rect 1726 28843 1782 28899
rect 1850 28843 1906 28899
rect 114 28719 170 28775
rect 238 28719 294 28775
rect 362 28719 418 28775
rect 486 28719 542 28775
rect 610 28719 666 28775
rect 734 28719 790 28775
rect 858 28719 914 28775
rect 982 28719 1038 28775
rect 1106 28719 1162 28775
rect 1230 28719 1286 28775
rect 1354 28719 1410 28775
rect 1478 28719 1534 28775
rect 1602 28719 1658 28775
rect 1726 28719 1782 28775
rect 1850 28719 1906 28775
rect 114 28595 170 28651
rect 238 28595 294 28651
rect 362 28595 418 28651
rect 486 28595 542 28651
rect 610 28595 666 28651
rect 734 28595 790 28651
rect 858 28595 914 28651
rect 982 28595 1038 28651
rect 1106 28595 1162 28651
rect 1230 28595 1286 28651
rect 1354 28595 1410 28651
rect 1478 28595 1534 28651
rect 1602 28595 1658 28651
rect 1726 28595 1782 28651
rect 1850 28595 1906 28651
rect 114 28471 170 28527
rect 238 28471 294 28527
rect 362 28471 418 28527
rect 486 28471 542 28527
rect 610 28471 666 28527
rect 734 28471 790 28527
rect 858 28471 914 28527
rect 982 28471 1038 28527
rect 1106 28471 1162 28527
rect 1230 28471 1286 28527
rect 1354 28471 1410 28527
rect 1478 28471 1534 28527
rect 1602 28471 1658 28527
rect 1726 28471 1782 28527
rect 1850 28471 1906 28527
rect 114 28347 170 28403
rect 238 28347 294 28403
rect 362 28347 418 28403
rect 486 28347 542 28403
rect 610 28347 666 28403
rect 734 28347 790 28403
rect 858 28347 914 28403
rect 982 28347 1038 28403
rect 1106 28347 1162 28403
rect 1230 28347 1286 28403
rect 1354 28347 1410 28403
rect 1478 28347 1534 28403
rect 1602 28347 1658 28403
rect 1726 28347 1782 28403
rect 1850 28347 1906 28403
rect 114 28223 170 28279
rect 238 28223 294 28279
rect 362 28223 418 28279
rect 486 28223 542 28279
rect 610 28223 666 28279
rect 734 28223 790 28279
rect 858 28223 914 28279
rect 982 28223 1038 28279
rect 1106 28223 1162 28279
rect 1230 28223 1286 28279
rect 1354 28223 1410 28279
rect 1478 28223 1534 28279
rect 1602 28223 1658 28279
rect 1726 28223 1782 28279
rect 1850 28223 1906 28279
rect 114 28099 170 28155
rect 238 28099 294 28155
rect 362 28099 418 28155
rect 486 28099 542 28155
rect 610 28099 666 28155
rect 734 28099 790 28155
rect 858 28099 914 28155
rect 982 28099 1038 28155
rect 1106 28099 1162 28155
rect 1230 28099 1286 28155
rect 1354 28099 1410 28155
rect 1478 28099 1534 28155
rect 1602 28099 1658 28155
rect 1726 28099 1782 28155
rect 1850 28099 1906 28155
rect 114 27975 170 28031
rect 238 27975 294 28031
rect 362 27975 418 28031
rect 486 27975 542 28031
rect 610 27975 666 28031
rect 734 27975 790 28031
rect 858 27975 914 28031
rect 982 27975 1038 28031
rect 1106 27975 1162 28031
rect 1230 27975 1286 28031
rect 1354 27975 1410 28031
rect 1478 27975 1534 28031
rect 1602 27975 1658 28031
rect 1726 27975 1782 28031
rect 1850 27975 1906 28031
rect 114 27851 170 27907
rect 238 27851 294 27907
rect 362 27851 418 27907
rect 486 27851 542 27907
rect 610 27851 666 27907
rect 734 27851 790 27907
rect 858 27851 914 27907
rect 982 27851 1038 27907
rect 1106 27851 1162 27907
rect 1230 27851 1286 27907
rect 1354 27851 1410 27907
rect 1478 27851 1534 27907
rect 1602 27851 1658 27907
rect 1726 27851 1782 27907
rect 1850 27851 1906 27907
rect 114 27727 170 27783
rect 238 27727 294 27783
rect 362 27727 418 27783
rect 486 27727 542 27783
rect 610 27727 666 27783
rect 734 27727 790 27783
rect 858 27727 914 27783
rect 982 27727 1038 27783
rect 1106 27727 1162 27783
rect 1230 27727 1286 27783
rect 1354 27727 1410 27783
rect 1478 27727 1534 27783
rect 1602 27727 1658 27783
rect 1726 27727 1782 27783
rect 1850 27727 1906 27783
rect 114 27603 170 27659
rect 238 27603 294 27659
rect 362 27603 418 27659
rect 486 27603 542 27659
rect 610 27603 666 27659
rect 734 27603 790 27659
rect 858 27603 914 27659
rect 982 27603 1038 27659
rect 1106 27603 1162 27659
rect 1230 27603 1286 27659
rect 1354 27603 1410 27659
rect 1478 27603 1534 27659
rect 1602 27603 1658 27659
rect 1726 27603 1782 27659
rect 1850 27603 1906 27659
rect 114 27479 170 27535
rect 238 27479 294 27535
rect 362 27479 418 27535
rect 486 27479 542 27535
rect 610 27479 666 27535
rect 734 27479 790 27535
rect 858 27479 914 27535
rect 982 27479 1038 27535
rect 1106 27479 1162 27535
rect 1230 27479 1286 27535
rect 1354 27479 1410 27535
rect 1478 27479 1534 27535
rect 1602 27479 1658 27535
rect 1726 27479 1782 27535
rect 1850 27479 1906 27535
rect 114 27355 170 27411
rect 238 27355 294 27411
rect 362 27355 418 27411
rect 486 27355 542 27411
rect 610 27355 666 27411
rect 734 27355 790 27411
rect 858 27355 914 27411
rect 982 27355 1038 27411
rect 1106 27355 1162 27411
rect 1230 27355 1286 27411
rect 1354 27355 1410 27411
rect 1478 27355 1534 27411
rect 1602 27355 1658 27411
rect 1726 27355 1782 27411
rect 1850 27355 1906 27411
rect 114 27231 170 27287
rect 238 27231 294 27287
rect 362 27231 418 27287
rect 486 27231 542 27287
rect 610 27231 666 27287
rect 734 27231 790 27287
rect 858 27231 914 27287
rect 982 27231 1038 27287
rect 1106 27231 1162 27287
rect 1230 27231 1286 27287
rect 1354 27231 1410 27287
rect 1478 27231 1534 27287
rect 1602 27231 1658 27287
rect 1726 27231 1782 27287
rect 1850 27231 1906 27287
rect 114 27107 170 27163
rect 238 27107 294 27163
rect 362 27107 418 27163
rect 486 27107 542 27163
rect 610 27107 666 27163
rect 734 27107 790 27163
rect 858 27107 914 27163
rect 982 27107 1038 27163
rect 1106 27107 1162 27163
rect 1230 27107 1286 27163
rect 1354 27107 1410 27163
rect 1478 27107 1534 27163
rect 1602 27107 1658 27163
rect 1726 27107 1782 27163
rect 1850 27107 1906 27163
rect 114 26983 170 27039
rect 238 26983 294 27039
rect 362 26983 418 27039
rect 486 26983 542 27039
rect 610 26983 666 27039
rect 734 26983 790 27039
rect 858 26983 914 27039
rect 982 26983 1038 27039
rect 1106 26983 1162 27039
rect 1230 26983 1286 27039
rect 1354 26983 1410 27039
rect 1478 26983 1534 27039
rect 1602 26983 1658 27039
rect 1726 26983 1782 27039
rect 1850 26983 1906 27039
rect 114 26445 170 26501
rect 238 26445 294 26501
rect 362 26445 418 26501
rect 486 26445 542 26501
rect 610 26445 666 26501
rect 734 26445 790 26501
rect 858 26445 914 26501
rect 982 26445 1038 26501
rect 1106 26445 1162 26501
rect 1230 26445 1286 26501
rect 1354 26445 1410 26501
rect 1478 26445 1534 26501
rect 1602 26445 1658 26501
rect 1726 26445 1782 26501
rect 1850 26445 1906 26501
rect 114 26321 170 26377
rect 238 26321 294 26377
rect 362 26321 418 26377
rect 486 26321 542 26377
rect 610 26321 666 26377
rect 734 26321 790 26377
rect 858 26321 914 26377
rect 982 26321 1038 26377
rect 1106 26321 1162 26377
rect 1230 26321 1286 26377
rect 1354 26321 1410 26377
rect 1478 26321 1534 26377
rect 1602 26321 1658 26377
rect 1726 26321 1782 26377
rect 1850 26321 1906 26377
rect 114 26197 170 26253
rect 238 26197 294 26253
rect 362 26197 418 26253
rect 486 26197 542 26253
rect 610 26197 666 26253
rect 734 26197 790 26253
rect 858 26197 914 26253
rect 982 26197 1038 26253
rect 1106 26197 1162 26253
rect 1230 26197 1286 26253
rect 1354 26197 1410 26253
rect 1478 26197 1534 26253
rect 1602 26197 1658 26253
rect 1726 26197 1782 26253
rect 1850 26197 1906 26253
rect 114 26073 170 26129
rect 238 26073 294 26129
rect 362 26073 418 26129
rect 486 26073 542 26129
rect 610 26073 666 26129
rect 734 26073 790 26129
rect 858 26073 914 26129
rect 982 26073 1038 26129
rect 1106 26073 1162 26129
rect 1230 26073 1286 26129
rect 1354 26073 1410 26129
rect 1478 26073 1534 26129
rect 1602 26073 1658 26129
rect 1726 26073 1782 26129
rect 1850 26073 1906 26129
rect 114 25949 170 26005
rect 238 25949 294 26005
rect 362 25949 418 26005
rect 486 25949 542 26005
rect 610 25949 666 26005
rect 734 25949 790 26005
rect 858 25949 914 26005
rect 982 25949 1038 26005
rect 1106 25949 1162 26005
rect 1230 25949 1286 26005
rect 1354 25949 1410 26005
rect 1478 25949 1534 26005
rect 1602 25949 1658 26005
rect 1726 25949 1782 26005
rect 1850 25949 1906 26005
rect 114 25825 170 25881
rect 238 25825 294 25881
rect 362 25825 418 25881
rect 486 25825 542 25881
rect 610 25825 666 25881
rect 734 25825 790 25881
rect 858 25825 914 25881
rect 982 25825 1038 25881
rect 1106 25825 1162 25881
rect 1230 25825 1286 25881
rect 1354 25825 1410 25881
rect 1478 25825 1534 25881
rect 1602 25825 1658 25881
rect 1726 25825 1782 25881
rect 1850 25825 1906 25881
rect 114 25701 170 25757
rect 238 25701 294 25757
rect 362 25701 418 25757
rect 486 25701 542 25757
rect 610 25701 666 25757
rect 734 25701 790 25757
rect 858 25701 914 25757
rect 982 25701 1038 25757
rect 1106 25701 1162 25757
rect 1230 25701 1286 25757
rect 1354 25701 1410 25757
rect 1478 25701 1534 25757
rect 1602 25701 1658 25757
rect 1726 25701 1782 25757
rect 1850 25701 1906 25757
rect 114 25577 170 25633
rect 238 25577 294 25633
rect 362 25577 418 25633
rect 486 25577 542 25633
rect 610 25577 666 25633
rect 734 25577 790 25633
rect 858 25577 914 25633
rect 982 25577 1038 25633
rect 1106 25577 1162 25633
rect 1230 25577 1286 25633
rect 1354 25577 1410 25633
rect 1478 25577 1534 25633
rect 1602 25577 1658 25633
rect 1726 25577 1782 25633
rect 1850 25577 1906 25633
rect 114 25453 170 25509
rect 238 25453 294 25509
rect 362 25453 418 25509
rect 486 25453 542 25509
rect 610 25453 666 25509
rect 734 25453 790 25509
rect 858 25453 914 25509
rect 982 25453 1038 25509
rect 1106 25453 1162 25509
rect 1230 25453 1286 25509
rect 1354 25453 1410 25509
rect 1478 25453 1534 25509
rect 1602 25453 1658 25509
rect 1726 25453 1782 25509
rect 1850 25453 1906 25509
rect 114 25329 170 25385
rect 238 25329 294 25385
rect 362 25329 418 25385
rect 486 25329 542 25385
rect 610 25329 666 25385
rect 734 25329 790 25385
rect 858 25329 914 25385
rect 982 25329 1038 25385
rect 1106 25329 1162 25385
rect 1230 25329 1286 25385
rect 1354 25329 1410 25385
rect 1478 25329 1534 25385
rect 1602 25329 1658 25385
rect 1726 25329 1782 25385
rect 1850 25329 1906 25385
rect 114 24832 170 24888
rect 238 24832 294 24888
rect 362 24832 418 24888
rect 486 24832 542 24888
rect 610 24832 666 24888
rect 734 24832 790 24888
rect 858 24832 914 24888
rect 982 24832 1038 24888
rect 1106 24832 1162 24888
rect 1230 24832 1286 24888
rect 1354 24832 1410 24888
rect 1478 24832 1534 24888
rect 1602 24832 1658 24888
rect 1726 24832 1782 24888
rect 1850 24832 1906 24888
rect 114 24708 170 24764
rect 238 24708 294 24764
rect 362 24708 418 24764
rect 486 24708 542 24764
rect 610 24708 666 24764
rect 734 24708 790 24764
rect 858 24708 914 24764
rect 982 24708 1038 24764
rect 1106 24708 1162 24764
rect 1230 24708 1286 24764
rect 1354 24708 1410 24764
rect 1478 24708 1534 24764
rect 1602 24708 1658 24764
rect 1726 24708 1782 24764
rect 1850 24708 1906 24764
rect 114 24584 170 24640
rect 238 24584 294 24640
rect 362 24584 418 24640
rect 486 24584 542 24640
rect 610 24584 666 24640
rect 734 24584 790 24640
rect 858 24584 914 24640
rect 982 24584 1038 24640
rect 1106 24584 1162 24640
rect 1230 24584 1286 24640
rect 1354 24584 1410 24640
rect 1478 24584 1534 24640
rect 1602 24584 1658 24640
rect 1726 24584 1782 24640
rect 1850 24584 1906 24640
rect 114 24460 170 24516
rect 238 24460 294 24516
rect 362 24460 418 24516
rect 486 24460 542 24516
rect 610 24460 666 24516
rect 734 24460 790 24516
rect 858 24460 914 24516
rect 982 24460 1038 24516
rect 1106 24460 1162 24516
rect 1230 24460 1286 24516
rect 1354 24460 1410 24516
rect 1478 24460 1534 24516
rect 1602 24460 1658 24516
rect 1726 24460 1782 24516
rect 1850 24460 1906 24516
rect 114 24336 170 24392
rect 238 24336 294 24392
rect 362 24336 418 24392
rect 486 24336 542 24392
rect 610 24336 666 24392
rect 734 24336 790 24392
rect 858 24336 914 24392
rect 982 24336 1038 24392
rect 1106 24336 1162 24392
rect 1230 24336 1286 24392
rect 1354 24336 1410 24392
rect 1478 24336 1534 24392
rect 1602 24336 1658 24392
rect 1726 24336 1782 24392
rect 1850 24336 1906 24392
rect 114 24212 170 24268
rect 238 24212 294 24268
rect 362 24212 418 24268
rect 486 24212 542 24268
rect 610 24212 666 24268
rect 734 24212 790 24268
rect 858 24212 914 24268
rect 982 24212 1038 24268
rect 1106 24212 1162 24268
rect 1230 24212 1286 24268
rect 1354 24212 1410 24268
rect 1478 24212 1534 24268
rect 1602 24212 1658 24268
rect 1726 24212 1782 24268
rect 1850 24212 1906 24268
rect 114 24088 170 24144
rect 238 24088 294 24144
rect 362 24088 418 24144
rect 486 24088 542 24144
rect 610 24088 666 24144
rect 734 24088 790 24144
rect 858 24088 914 24144
rect 982 24088 1038 24144
rect 1106 24088 1162 24144
rect 1230 24088 1286 24144
rect 1354 24088 1410 24144
rect 1478 24088 1534 24144
rect 1602 24088 1658 24144
rect 1726 24088 1782 24144
rect 1850 24088 1906 24144
rect 114 23964 170 24020
rect 238 23964 294 24020
rect 362 23964 418 24020
rect 486 23964 542 24020
rect 610 23964 666 24020
rect 734 23964 790 24020
rect 858 23964 914 24020
rect 982 23964 1038 24020
rect 1106 23964 1162 24020
rect 1230 23964 1286 24020
rect 1354 23964 1410 24020
rect 1478 23964 1534 24020
rect 1602 23964 1658 24020
rect 1726 23964 1782 24020
rect 1850 23964 1906 24020
rect 114 23840 170 23896
rect 238 23840 294 23896
rect 362 23840 418 23896
rect 486 23840 542 23896
rect 610 23840 666 23896
rect 734 23840 790 23896
rect 858 23840 914 23896
rect 982 23840 1038 23896
rect 1106 23840 1162 23896
rect 1230 23840 1286 23896
rect 1354 23840 1410 23896
rect 1478 23840 1534 23896
rect 1602 23840 1658 23896
rect 1726 23840 1782 23896
rect 1850 23840 1906 23896
rect 114 23716 170 23772
rect 238 23716 294 23772
rect 362 23716 418 23772
rect 486 23716 542 23772
rect 610 23716 666 23772
rect 734 23716 790 23772
rect 858 23716 914 23772
rect 982 23716 1038 23772
rect 1106 23716 1162 23772
rect 1230 23716 1286 23772
rect 1354 23716 1410 23772
rect 1478 23716 1534 23772
rect 1602 23716 1658 23772
rect 1726 23716 1782 23772
rect 1850 23716 1906 23772
rect 114 23178 170 23234
rect 238 23178 294 23234
rect 362 23178 418 23234
rect 486 23178 542 23234
rect 610 23178 666 23234
rect 734 23178 790 23234
rect 858 23178 914 23234
rect 982 23178 1038 23234
rect 1106 23178 1162 23234
rect 1230 23178 1286 23234
rect 1354 23178 1410 23234
rect 1478 23178 1534 23234
rect 1602 23178 1658 23234
rect 1726 23178 1782 23234
rect 1850 23178 1906 23234
rect 114 23054 170 23110
rect 238 23054 294 23110
rect 362 23054 418 23110
rect 486 23054 542 23110
rect 610 23054 666 23110
rect 734 23054 790 23110
rect 858 23054 914 23110
rect 982 23054 1038 23110
rect 1106 23054 1162 23110
rect 1230 23054 1286 23110
rect 1354 23054 1410 23110
rect 1478 23054 1534 23110
rect 1602 23054 1658 23110
rect 1726 23054 1782 23110
rect 1850 23054 1906 23110
rect 114 22930 170 22986
rect 238 22930 294 22986
rect 362 22930 418 22986
rect 486 22930 542 22986
rect 610 22930 666 22986
rect 734 22930 790 22986
rect 858 22930 914 22986
rect 982 22930 1038 22986
rect 1106 22930 1162 22986
rect 1230 22930 1286 22986
rect 1354 22930 1410 22986
rect 1478 22930 1534 22986
rect 1602 22930 1658 22986
rect 1726 22930 1782 22986
rect 1850 22930 1906 22986
rect 114 22806 170 22862
rect 238 22806 294 22862
rect 362 22806 418 22862
rect 486 22806 542 22862
rect 610 22806 666 22862
rect 734 22806 790 22862
rect 858 22806 914 22862
rect 982 22806 1038 22862
rect 1106 22806 1162 22862
rect 1230 22806 1286 22862
rect 1354 22806 1410 22862
rect 1478 22806 1534 22862
rect 1602 22806 1658 22862
rect 1726 22806 1782 22862
rect 1850 22806 1906 22862
rect 114 22682 170 22738
rect 238 22682 294 22738
rect 362 22682 418 22738
rect 486 22682 542 22738
rect 610 22682 666 22738
rect 734 22682 790 22738
rect 858 22682 914 22738
rect 982 22682 1038 22738
rect 1106 22682 1162 22738
rect 1230 22682 1286 22738
rect 1354 22682 1410 22738
rect 1478 22682 1534 22738
rect 1602 22682 1658 22738
rect 1726 22682 1782 22738
rect 1850 22682 1906 22738
rect 114 22558 170 22614
rect 238 22558 294 22614
rect 362 22558 418 22614
rect 486 22558 542 22614
rect 610 22558 666 22614
rect 734 22558 790 22614
rect 858 22558 914 22614
rect 982 22558 1038 22614
rect 1106 22558 1162 22614
rect 1230 22558 1286 22614
rect 1354 22558 1410 22614
rect 1478 22558 1534 22614
rect 1602 22558 1658 22614
rect 1726 22558 1782 22614
rect 1850 22558 1906 22614
rect 114 22434 170 22490
rect 238 22434 294 22490
rect 362 22434 418 22490
rect 486 22434 542 22490
rect 610 22434 666 22490
rect 734 22434 790 22490
rect 858 22434 914 22490
rect 982 22434 1038 22490
rect 1106 22434 1162 22490
rect 1230 22434 1286 22490
rect 1354 22434 1410 22490
rect 1478 22434 1534 22490
rect 1602 22434 1658 22490
rect 1726 22434 1782 22490
rect 1850 22434 1906 22490
rect 114 22310 170 22366
rect 238 22310 294 22366
rect 362 22310 418 22366
rect 486 22310 542 22366
rect 610 22310 666 22366
rect 734 22310 790 22366
rect 858 22310 914 22366
rect 982 22310 1038 22366
rect 1106 22310 1162 22366
rect 1230 22310 1286 22366
rect 1354 22310 1410 22366
rect 1478 22310 1534 22366
rect 1602 22310 1658 22366
rect 1726 22310 1782 22366
rect 1850 22310 1906 22366
rect 114 22186 170 22242
rect 238 22186 294 22242
rect 362 22186 418 22242
rect 486 22186 542 22242
rect 610 22186 666 22242
rect 734 22186 790 22242
rect 858 22186 914 22242
rect 982 22186 1038 22242
rect 1106 22186 1162 22242
rect 1230 22186 1286 22242
rect 1354 22186 1410 22242
rect 1478 22186 1534 22242
rect 1602 22186 1658 22242
rect 1726 22186 1782 22242
rect 1850 22186 1906 22242
rect 114 22062 170 22118
rect 238 22062 294 22118
rect 362 22062 418 22118
rect 486 22062 542 22118
rect 610 22062 666 22118
rect 734 22062 790 22118
rect 858 22062 914 22118
rect 982 22062 1038 22118
rect 1106 22062 1162 22118
rect 1230 22062 1286 22118
rect 1354 22062 1410 22118
rect 1478 22062 1534 22118
rect 1602 22062 1658 22118
rect 1726 22062 1782 22118
rect 1850 22062 1906 22118
rect 114 21938 170 21994
rect 238 21938 294 21994
rect 362 21938 418 21994
rect 486 21938 542 21994
rect 610 21938 666 21994
rect 734 21938 790 21994
rect 858 21938 914 21994
rect 982 21938 1038 21994
rect 1106 21938 1162 21994
rect 1230 21938 1286 21994
rect 1354 21938 1410 21994
rect 1478 21938 1534 21994
rect 1602 21938 1658 21994
rect 1726 21938 1782 21994
rect 1850 21938 1906 21994
rect 114 21814 170 21870
rect 238 21814 294 21870
rect 362 21814 418 21870
rect 486 21814 542 21870
rect 610 21814 666 21870
rect 734 21814 790 21870
rect 858 21814 914 21870
rect 982 21814 1038 21870
rect 1106 21814 1162 21870
rect 1230 21814 1286 21870
rect 1354 21814 1410 21870
rect 1478 21814 1534 21870
rect 1602 21814 1658 21870
rect 1726 21814 1782 21870
rect 1850 21814 1906 21870
rect 114 21690 170 21746
rect 238 21690 294 21746
rect 362 21690 418 21746
rect 486 21690 542 21746
rect 610 21690 666 21746
rect 734 21690 790 21746
rect 858 21690 914 21746
rect 982 21690 1038 21746
rect 1106 21690 1162 21746
rect 1230 21690 1286 21746
rect 1354 21690 1410 21746
rect 1478 21690 1534 21746
rect 1602 21690 1658 21746
rect 1726 21690 1782 21746
rect 1850 21690 1906 21746
rect 114 21566 170 21622
rect 238 21566 294 21622
rect 362 21566 418 21622
rect 486 21566 542 21622
rect 610 21566 666 21622
rect 734 21566 790 21622
rect 858 21566 914 21622
rect 982 21566 1038 21622
rect 1106 21566 1162 21622
rect 1230 21566 1286 21622
rect 1354 21566 1410 21622
rect 1478 21566 1534 21622
rect 1602 21566 1658 21622
rect 1726 21566 1782 21622
rect 1850 21566 1906 21622
rect 114 21442 170 21498
rect 238 21442 294 21498
rect 362 21442 418 21498
rect 486 21442 542 21498
rect 610 21442 666 21498
rect 734 21442 790 21498
rect 858 21442 914 21498
rect 982 21442 1038 21498
rect 1106 21442 1162 21498
rect 1230 21442 1286 21498
rect 1354 21442 1410 21498
rect 1478 21442 1534 21498
rect 1602 21442 1658 21498
rect 1726 21442 1782 21498
rect 1850 21442 1906 21498
rect 114 21318 170 21374
rect 238 21318 294 21374
rect 362 21318 418 21374
rect 486 21318 542 21374
rect 610 21318 666 21374
rect 734 21318 790 21374
rect 858 21318 914 21374
rect 982 21318 1038 21374
rect 1106 21318 1162 21374
rect 1230 21318 1286 21374
rect 1354 21318 1410 21374
rect 1478 21318 1534 21374
rect 1602 21318 1658 21374
rect 1726 21318 1782 21374
rect 1850 21318 1906 21374
rect 114 21194 170 21250
rect 238 21194 294 21250
rect 362 21194 418 21250
rect 486 21194 542 21250
rect 610 21194 666 21250
rect 734 21194 790 21250
rect 858 21194 914 21250
rect 982 21194 1038 21250
rect 1106 21194 1162 21250
rect 1230 21194 1286 21250
rect 1354 21194 1410 21250
rect 1478 21194 1534 21250
rect 1602 21194 1658 21250
rect 1726 21194 1782 21250
rect 1850 21194 1906 21250
rect 114 21070 170 21126
rect 238 21070 294 21126
rect 362 21070 418 21126
rect 486 21070 542 21126
rect 610 21070 666 21126
rect 734 21070 790 21126
rect 858 21070 914 21126
rect 982 21070 1038 21126
rect 1106 21070 1162 21126
rect 1230 21070 1286 21126
rect 1354 21070 1410 21126
rect 1478 21070 1534 21126
rect 1602 21070 1658 21126
rect 1726 21070 1782 21126
rect 1850 21070 1906 21126
rect 114 20946 170 21002
rect 238 20946 294 21002
rect 362 20946 418 21002
rect 486 20946 542 21002
rect 610 20946 666 21002
rect 734 20946 790 21002
rect 858 20946 914 21002
rect 982 20946 1038 21002
rect 1106 20946 1162 21002
rect 1230 20946 1286 21002
rect 1354 20946 1410 21002
rect 1478 20946 1534 21002
rect 1602 20946 1658 21002
rect 1726 20946 1782 21002
rect 1850 20946 1906 21002
rect 114 20822 170 20878
rect 238 20822 294 20878
rect 362 20822 418 20878
rect 486 20822 542 20878
rect 610 20822 666 20878
rect 734 20822 790 20878
rect 858 20822 914 20878
rect 982 20822 1038 20878
rect 1106 20822 1162 20878
rect 1230 20822 1286 20878
rect 1354 20822 1410 20878
rect 1478 20822 1534 20878
rect 1602 20822 1658 20878
rect 1726 20822 1782 20878
rect 1850 20822 1906 20878
rect 114 20698 170 20754
rect 238 20698 294 20754
rect 362 20698 418 20754
rect 486 20698 542 20754
rect 610 20698 666 20754
rect 734 20698 790 20754
rect 858 20698 914 20754
rect 982 20698 1038 20754
rect 1106 20698 1162 20754
rect 1230 20698 1286 20754
rect 1354 20698 1410 20754
rect 1478 20698 1534 20754
rect 1602 20698 1658 20754
rect 1726 20698 1782 20754
rect 1850 20698 1906 20754
rect 114 20574 170 20630
rect 238 20574 294 20630
rect 362 20574 418 20630
rect 486 20574 542 20630
rect 610 20574 666 20630
rect 734 20574 790 20630
rect 858 20574 914 20630
rect 982 20574 1038 20630
rect 1106 20574 1162 20630
rect 1230 20574 1286 20630
rect 1354 20574 1410 20630
rect 1478 20574 1534 20630
rect 1602 20574 1658 20630
rect 1726 20574 1782 20630
rect 1850 20574 1906 20630
rect 114 19967 170 20023
rect 238 19967 294 20023
rect 362 19967 418 20023
rect 486 19967 542 20023
rect 610 19967 666 20023
rect 734 19967 790 20023
rect 858 19967 914 20023
rect 982 19967 1038 20023
rect 1106 19967 1162 20023
rect 1230 19967 1286 20023
rect 1354 19967 1410 20023
rect 1478 19967 1534 20023
rect 1602 19967 1658 20023
rect 1726 19967 1782 20023
rect 1850 19967 1906 20023
rect 114 19843 170 19899
rect 238 19843 294 19899
rect 362 19843 418 19899
rect 486 19843 542 19899
rect 610 19843 666 19899
rect 734 19843 790 19899
rect 858 19843 914 19899
rect 982 19843 1038 19899
rect 1106 19843 1162 19899
rect 1230 19843 1286 19899
rect 1354 19843 1410 19899
rect 1478 19843 1534 19899
rect 1602 19843 1658 19899
rect 1726 19843 1782 19899
rect 1850 19843 1906 19899
rect 114 19719 170 19775
rect 238 19719 294 19775
rect 362 19719 418 19775
rect 486 19719 542 19775
rect 610 19719 666 19775
rect 734 19719 790 19775
rect 858 19719 914 19775
rect 982 19719 1038 19775
rect 1106 19719 1162 19775
rect 1230 19719 1286 19775
rect 1354 19719 1410 19775
rect 1478 19719 1534 19775
rect 1602 19719 1658 19775
rect 1726 19719 1782 19775
rect 1850 19719 1906 19775
rect 114 19595 170 19651
rect 238 19595 294 19651
rect 362 19595 418 19651
rect 486 19595 542 19651
rect 610 19595 666 19651
rect 734 19595 790 19651
rect 858 19595 914 19651
rect 982 19595 1038 19651
rect 1106 19595 1162 19651
rect 1230 19595 1286 19651
rect 1354 19595 1410 19651
rect 1478 19595 1534 19651
rect 1602 19595 1658 19651
rect 1726 19595 1782 19651
rect 1850 19595 1906 19651
rect 114 19471 170 19527
rect 238 19471 294 19527
rect 362 19471 418 19527
rect 486 19471 542 19527
rect 610 19471 666 19527
rect 734 19471 790 19527
rect 858 19471 914 19527
rect 982 19471 1038 19527
rect 1106 19471 1162 19527
rect 1230 19471 1286 19527
rect 1354 19471 1410 19527
rect 1478 19471 1534 19527
rect 1602 19471 1658 19527
rect 1726 19471 1782 19527
rect 1850 19471 1906 19527
rect 114 19347 170 19403
rect 238 19347 294 19403
rect 362 19347 418 19403
rect 486 19347 542 19403
rect 610 19347 666 19403
rect 734 19347 790 19403
rect 858 19347 914 19403
rect 982 19347 1038 19403
rect 1106 19347 1162 19403
rect 1230 19347 1286 19403
rect 1354 19347 1410 19403
rect 1478 19347 1534 19403
rect 1602 19347 1658 19403
rect 1726 19347 1782 19403
rect 1850 19347 1906 19403
rect 114 19223 170 19279
rect 238 19223 294 19279
rect 362 19223 418 19279
rect 486 19223 542 19279
rect 610 19223 666 19279
rect 734 19223 790 19279
rect 858 19223 914 19279
rect 982 19223 1038 19279
rect 1106 19223 1162 19279
rect 1230 19223 1286 19279
rect 1354 19223 1410 19279
rect 1478 19223 1534 19279
rect 1602 19223 1658 19279
rect 1726 19223 1782 19279
rect 1850 19223 1906 19279
rect 114 19099 170 19155
rect 238 19099 294 19155
rect 362 19099 418 19155
rect 486 19099 542 19155
rect 610 19099 666 19155
rect 734 19099 790 19155
rect 858 19099 914 19155
rect 982 19099 1038 19155
rect 1106 19099 1162 19155
rect 1230 19099 1286 19155
rect 1354 19099 1410 19155
rect 1478 19099 1534 19155
rect 1602 19099 1658 19155
rect 1726 19099 1782 19155
rect 1850 19099 1906 19155
rect 114 18975 170 19031
rect 238 18975 294 19031
rect 362 18975 418 19031
rect 486 18975 542 19031
rect 610 18975 666 19031
rect 734 18975 790 19031
rect 858 18975 914 19031
rect 982 18975 1038 19031
rect 1106 18975 1162 19031
rect 1230 18975 1286 19031
rect 1354 18975 1410 19031
rect 1478 18975 1534 19031
rect 1602 18975 1658 19031
rect 1726 18975 1782 19031
rect 1850 18975 1906 19031
rect 114 18851 170 18907
rect 238 18851 294 18907
rect 362 18851 418 18907
rect 486 18851 542 18907
rect 610 18851 666 18907
rect 734 18851 790 18907
rect 858 18851 914 18907
rect 982 18851 1038 18907
rect 1106 18851 1162 18907
rect 1230 18851 1286 18907
rect 1354 18851 1410 18907
rect 1478 18851 1534 18907
rect 1602 18851 1658 18907
rect 1726 18851 1782 18907
rect 1850 18851 1906 18907
rect 114 18727 170 18783
rect 238 18727 294 18783
rect 362 18727 418 18783
rect 486 18727 542 18783
rect 610 18727 666 18783
rect 734 18727 790 18783
rect 858 18727 914 18783
rect 982 18727 1038 18783
rect 1106 18727 1162 18783
rect 1230 18727 1286 18783
rect 1354 18727 1410 18783
rect 1478 18727 1534 18783
rect 1602 18727 1658 18783
rect 1726 18727 1782 18783
rect 1850 18727 1906 18783
rect 114 18603 170 18659
rect 238 18603 294 18659
rect 362 18603 418 18659
rect 486 18603 542 18659
rect 610 18603 666 18659
rect 734 18603 790 18659
rect 858 18603 914 18659
rect 982 18603 1038 18659
rect 1106 18603 1162 18659
rect 1230 18603 1286 18659
rect 1354 18603 1410 18659
rect 1478 18603 1534 18659
rect 1602 18603 1658 18659
rect 1726 18603 1782 18659
rect 1850 18603 1906 18659
rect 114 18479 170 18535
rect 238 18479 294 18535
rect 362 18479 418 18535
rect 486 18479 542 18535
rect 610 18479 666 18535
rect 734 18479 790 18535
rect 858 18479 914 18535
rect 982 18479 1038 18535
rect 1106 18479 1162 18535
rect 1230 18479 1286 18535
rect 1354 18479 1410 18535
rect 1478 18479 1534 18535
rect 1602 18479 1658 18535
rect 1726 18479 1782 18535
rect 1850 18479 1906 18535
rect 114 18355 170 18411
rect 238 18355 294 18411
rect 362 18355 418 18411
rect 486 18355 542 18411
rect 610 18355 666 18411
rect 734 18355 790 18411
rect 858 18355 914 18411
rect 982 18355 1038 18411
rect 1106 18355 1162 18411
rect 1230 18355 1286 18411
rect 1354 18355 1410 18411
rect 1478 18355 1534 18411
rect 1602 18355 1658 18411
rect 1726 18355 1782 18411
rect 1850 18355 1906 18411
rect 114 18231 170 18287
rect 238 18231 294 18287
rect 362 18231 418 18287
rect 486 18231 542 18287
rect 610 18231 666 18287
rect 734 18231 790 18287
rect 858 18231 914 18287
rect 982 18231 1038 18287
rect 1106 18231 1162 18287
rect 1230 18231 1286 18287
rect 1354 18231 1410 18287
rect 1478 18231 1534 18287
rect 1602 18231 1658 18287
rect 1726 18231 1782 18287
rect 1850 18231 1906 18287
rect 114 18107 170 18163
rect 238 18107 294 18163
rect 362 18107 418 18163
rect 486 18107 542 18163
rect 610 18107 666 18163
rect 734 18107 790 18163
rect 858 18107 914 18163
rect 982 18107 1038 18163
rect 1106 18107 1162 18163
rect 1230 18107 1286 18163
rect 1354 18107 1410 18163
rect 1478 18107 1534 18163
rect 1602 18107 1658 18163
rect 1726 18107 1782 18163
rect 1850 18107 1906 18163
rect 114 17983 170 18039
rect 238 17983 294 18039
rect 362 17983 418 18039
rect 486 17983 542 18039
rect 610 17983 666 18039
rect 734 17983 790 18039
rect 858 17983 914 18039
rect 982 17983 1038 18039
rect 1106 17983 1162 18039
rect 1230 17983 1286 18039
rect 1354 17983 1410 18039
rect 1478 17983 1534 18039
rect 1602 17983 1658 18039
rect 1726 17983 1782 18039
rect 1850 17983 1906 18039
rect 114 17859 170 17915
rect 238 17859 294 17915
rect 362 17859 418 17915
rect 486 17859 542 17915
rect 610 17859 666 17915
rect 734 17859 790 17915
rect 858 17859 914 17915
rect 982 17859 1038 17915
rect 1106 17859 1162 17915
rect 1230 17859 1286 17915
rect 1354 17859 1410 17915
rect 1478 17859 1534 17915
rect 1602 17859 1658 17915
rect 1726 17859 1782 17915
rect 1850 17859 1906 17915
rect 114 17735 170 17791
rect 238 17735 294 17791
rect 362 17735 418 17791
rect 486 17735 542 17791
rect 610 17735 666 17791
rect 734 17735 790 17791
rect 858 17735 914 17791
rect 982 17735 1038 17791
rect 1106 17735 1162 17791
rect 1230 17735 1286 17791
rect 1354 17735 1410 17791
rect 1478 17735 1534 17791
rect 1602 17735 1658 17791
rect 1726 17735 1782 17791
rect 1850 17735 1906 17791
rect 114 17611 170 17667
rect 238 17611 294 17667
rect 362 17611 418 17667
rect 486 17611 542 17667
rect 610 17611 666 17667
rect 734 17611 790 17667
rect 858 17611 914 17667
rect 982 17611 1038 17667
rect 1106 17611 1162 17667
rect 1230 17611 1286 17667
rect 1354 17611 1410 17667
rect 1478 17611 1534 17667
rect 1602 17611 1658 17667
rect 1726 17611 1782 17667
rect 1850 17611 1906 17667
rect 114 17487 170 17543
rect 238 17487 294 17543
rect 362 17487 418 17543
rect 486 17487 542 17543
rect 610 17487 666 17543
rect 734 17487 790 17543
rect 858 17487 914 17543
rect 982 17487 1038 17543
rect 1106 17487 1162 17543
rect 1230 17487 1286 17543
rect 1354 17487 1410 17543
rect 1478 17487 1534 17543
rect 1602 17487 1658 17543
rect 1726 17487 1782 17543
rect 1850 17487 1906 17543
rect 114 17363 170 17419
rect 238 17363 294 17419
rect 362 17363 418 17419
rect 486 17363 542 17419
rect 610 17363 666 17419
rect 734 17363 790 17419
rect 858 17363 914 17419
rect 982 17363 1038 17419
rect 1106 17363 1162 17419
rect 1230 17363 1286 17419
rect 1354 17363 1410 17419
rect 1478 17363 1534 17419
rect 1602 17363 1658 17419
rect 1726 17363 1782 17419
rect 1850 17363 1906 17419
rect 114 16796 170 16852
rect 238 16796 294 16852
rect 362 16796 418 16852
rect 486 16796 542 16852
rect 610 16796 666 16852
rect 734 16796 790 16852
rect 858 16796 914 16852
rect 982 16796 1038 16852
rect 1106 16796 1162 16852
rect 1230 16796 1286 16852
rect 1354 16796 1410 16852
rect 1478 16796 1534 16852
rect 1602 16796 1658 16852
rect 1726 16796 1782 16852
rect 1850 16796 1906 16852
rect 114 16672 170 16728
rect 238 16672 294 16728
rect 362 16672 418 16728
rect 486 16672 542 16728
rect 610 16672 666 16728
rect 734 16672 790 16728
rect 858 16672 914 16728
rect 982 16672 1038 16728
rect 1106 16672 1162 16728
rect 1230 16672 1286 16728
rect 1354 16672 1410 16728
rect 1478 16672 1534 16728
rect 1602 16672 1658 16728
rect 1726 16672 1782 16728
rect 1850 16672 1906 16728
rect 114 16548 170 16604
rect 238 16548 294 16604
rect 362 16548 418 16604
rect 486 16548 542 16604
rect 610 16548 666 16604
rect 734 16548 790 16604
rect 858 16548 914 16604
rect 982 16548 1038 16604
rect 1106 16548 1162 16604
rect 1230 16548 1286 16604
rect 1354 16548 1410 16604
rect 1478 16548 1534 16604
rect 1602 16548 1658 16604
rect 1726 16548 1782 16604
rect 1850 16548 1906 16604
rect 114 16424 170 16480
rect 238 16424 294 16480
rect 362 16424 418 16480
rect 486 16424 542 16480
rect 610 16424 666 16480
rect 734 16424 790 16480
rect 858 16424 914 16480
rect 982 16424 1038 16480
rect 1106 16424 1162 16480
rect 1230 16424 1286 16480
rect 1354 16424 1410 16480
rect 1478 16424 1534 16480
rect 1602 16424 1658 16480
rect 1726 16424 1782 16480
rect 1850 16424 1906 16480
rect 114 16300 170 16356
rect 238 16300 294 16356
rect 362 16300 418 16356
rect 486 16300 542 16356
rect 610 16300 666 16356
rect 734 16300 790 16356
rect 858 16300 914 16356
rect 982 16300 1038 16356
rect 1106 16300 1162 16356
rect 1230 16300 1286 16356
rect 1354 16300 1410 16356
rect 1478 16300 1534 16356
rect 1602 16300 1658 16356
rect 1726 16300 1782 16356
rect 1850 16300 1906 16356
rect 114 16176 170 16232
rect 238 16176 294 16232
rect 362 16176 418 16232
rect 486 16176 542 16232
rect 610 16176 666 16232
rect 734 16176 790 16232
rect 858 16176 914 16232
rect 982 16176 1038 16232
rect 1106 16176 1162 16232
rect 1230 16176 1286 16232
rect 1354 16176 1410 16232
rect 1478 16176 1534 16232
rect 1602 16176 1658 16232
rect 1726 16176 1782 16232
rect 1850 16176 1906 16232
rect 114 16052 170 16108
rect 238 16052 294 16108
rect 362 16052 418 16108
rect 486 16052 542 16108
rect 610 16052 666 16108
rect 734 16052 790 16108
rect 858 16052 914 16108
rect 982 16052 1038 16108
rect 1106 16052 1162 16108
rect 1230 16052 1286 16108
rect 1354 16052 1410 16108
rect 1478 16052 1534 16108
rect 1602 16052 1658 16108
rect 1726 16052 1782 16108
rect 1850 16052 1906 16108
rect 114 15928 170 15984
rect 238 15928 294 15984
rect 362 15928 418 15984
rect 486 15928 542 15984
rect 610 15928 666 15984
rect 734 15928 790 15984
rect 858 15928 914 15984
rect 982 15928 1038 15984
rect 1106 15928 1162 15984
rect 1230 15928 1286 15984
rect 1354 15928 1410 15984
rect 1478 15928 1534 15984
rect 1602 15928 1658 15984
rect 1726 15928 1782 15984
rect 1850 15928 1906 15984
rect 114 15804 170 15860
rect 238 15804 294 15860
rect 362 15804 418 15860
rect 486 15804 542 15860
rect 610 15804 666 15860
rect 734 15804 790 15860
rect 858 15804 914 15860
rect 982 15804 1038 15860
rect 1106 15804 1162 15860
rect 1230 15804 1286 15860
rect 1354 15804 1410 15860
rect 1478 15804 1534 15860
rect 1602 15804 1658 15860
rect 1726 15804 1782 15860
rect 1850 15804 1906 15860
rect 114 15680 170 15736
rect 238 15680 294 15736
rect 362 15680 418 15736
rect 486 15680 542 15736
rect 610 15680 666 15736
rect 734 15680 790 15736
rect 858 15680 914 15736
rect 982 15680 1038 15736
rect 1106 15680 1162 15736
rect 1230 15680 1286 15736
rect 1354 15680 1410 15736
rect 1478 15680 1534 15736
rect 1602 15680 1658 15736
rect 1726 15680 1782 15736
rect 1850 15680 1906 15736
rect 114 15556 170 15612
rect 238 15556 294 15612
rect 362 15556 418 15612
rect 486 15556 542 15612
rect 610 15556 666 15612
rect 734 15556 790 15612
rect 858 15556 914 15612
rect 982 15556 1038 15612
rect 1106 15556 1162 15612
rect 1230 15556 1286 15612
rect 1354 15556 1410 15612
rect 1478 15556 1534 15612
rect 1602 15556 1658 15612
rect 1726 15556 1782 15612
rect 1850 15556 1906 15612
rect 114 15432 170 15488
rect 238 15432 294 15488
rect 362 15432 418 15488
rect 486 15432 542 15488
rect 610 15432 666 15488
rect 734 15432 790 15488
rect 858 15432 914 15488
rect 982 15432 1038 15488
rect 1106 15432 1162 15488
rect 1230 15432 1286 15488
rect 1354 15432 1410 15488
rect 1478 15432 1534 15488
rect 1602 15432 1658 15488
rect 1726 15432 1782 15488
rect 1850 15432 1906 15488
rect 114 15308 170 15364
rect 238 15308 294 15364
rect 362 15308 418 15364
rect 486 15308 542 15364
rect 610 15308 666 15364
rect 734 15308 790 15364
rect 858 15308 914 15364
rect 982 15308 1038 15364
rect 1106 15308 1162 15364
rect 1230 15308 1286 15364
rect 1354 15308 1410 15364
rect 1478 15308 1534 15364
rect 1602 15308 1658 15364
rect 1726 15308 1782 15364
rect 1850 15308 1906 15364
rect 114 15184 170 15240
rect 238 15184 294 15240
rect 362 15184 418 15240
rect 486 15184 542 15240
rect 610 15184 666 15240
rect 734 15184 790 15240
rect 858 15184 914 15240
rect 982 15184 1038 15240
rect 1106 15184 1162 15240
rect 1230 15184 1286 15240
rect 1354 15184 1410 15240
rect 1478 15184 1534 15240
rect 1602 15184 1658 15240
rect 1726 15184 1782 15240
rect 1850 15184 1906 15240
rect 114 15060 170 15116
rect 238 15060 294 15116
rect 362 15060 418 15116
rect 486 15060 542 15116
rect 610 15060 666 15116
rect 734 15060 790 15116
rect 858 15060 914 15116
rect 982 15060 1038 15116
rect 1106 15060 1162 15116
rect 1230 15060 1286 15116
rect 1354 15060 1410 15116
rect 1478 15060 1534 15116
rect 1602 15060 1658 15116
rect 1726 15060 1782 15116
rect 1850 15060 1906 15116
rect 114 14936 170 14992
rect 238 14936 294 14992
rect 362 14936 418 14992
rect 486 14936 542 14992
rect 610 14936 666 14992
rect 734 14936 790 14992
rect 858 14936 914 14992
rect 982 14936 1038 14992
rect 1106 14936 1162 14992
rect 1230 14936 1286 14992
rect 1354 14936 1410 14992
rect 1478 14936 1534 14992
rect 1602 14936 1658 14992
rect 1726 14936 1782 14992
rect 1850 14936 1906 14992
rect 114 14812 170 14868
rect 238 14812 294 14868
rect 362 14812 418 14868
rect 486 14812 542 14868
rect 610 14812 666 14868
rect 734 14812 790 14868
rect 858 14812 914 14868
rect 982 14812 1038 14868
rect 1106 14812 1162 14868
rect 1230 14812 1286 14868
rect 1354 14812 1410 14868
rect 1478 14812 1534 14868
rect 1602 14812 1658 14868
rect 1726 14812 1782 14868
rect 1850 14812 1906 14868
rect 114 14688 170 14744
rect 238 14688 294 14744
rect 362 14688 418 14744
rect 486 14688 542 14744
rect 610 14688 666 14744
rect 734 14688 790 14744
rect 858 14688 914 14744
rect 982 14688 1038 14744
rect 1106 14688 1162 14744
rect 1230 14688 1286 14744
rect 1354 14688 1410 14744
rect 1478 14688 1534 14744
rect 1602 14688 1658 14744
rect 1726 14688 1782 14744
rect 1850 14688 1906 14744
rect 114 14564 170 14620
rect 238 14564 294 14620
rect 362 14564 418 14620
rect 486 14564 542 14620
rect 610 14564 666 14620
rect 734 14564 790 14620
rect 858 14564 914 14620
rect 982 14564 1038 14620
rect 1106 14564 1162 14620
rect 1230 14564 1286 14620
rect 1354 14564 1410 14620
rect 1478 14564 1534 14620
rect 1602 14564 1658 14620
rect 1726 14564 1782 14620
rect 1850 14564 1906 14620
rect 114 14440 170 14496
rect 238 14440 294 14496
rect 362 14440 418 14496
rect 486 14440 542 14496
rect 610 14440 666 14496
rect 734 14440 790 14496
rect 858 14440 914 14496
rect 982 14440 1038 14496
rect 1106 14440 1162 14496
rect 1230 14440 1286 14496
rect 1354 14440 1410 14496
rect 1478 14440 1534 14496
rect 1602 14440 1658 14496
rect 1726 14440 1782 14496
rect 1850 14440 1906 14496
rect 114 14316 170 14372
rect 238 14316 294 14372
rect 362 14316 418 14372
rect 486 14316 542 14372
rect 610 14316 666 14372
rect 734 14316 790 14372
rect 858 14316 914 14372
rect 982 14316 1038 14372
rect 1106 14316 1162 14372
rect 1230 14316 1286 14372
rect 1354 14316 1410 14372
rect 1478 14316 1534 14372
rect 1602 14316 1658 14372
rect 1726 14316 1782 14372
rect 1850 14316 1906 14372
rect 114 14192 170 14248
rect 238 14192 294 14248
rect 362 14192 418 14248
rect 486 14192 542 14248
rect 610 14192 666 14248
rect 734 14192 790 14248
rect 858 14192 914 14248
rect 982 14192 1038 14248
rect 1106 14192 1162 14248
rect 1230 14192 1286 14248
rect 1354 14192 1410 14248
rect 1478 14192 1534 14248
rect 1602 14192 1658 14248
rect 1726 14192 1782 14248
rect 1850 14192 1906 14248
<< metal4 >>
rect 0 69624 2000 69678
rect 0 69568 114 69624
rect 170 69568 238 69624
rect 294 69568 362 69624
rect 418 69568 486 69624
rect 542 69568 610 69624
rect 666 69568 734 69624
rect 790 69568 858 69624
rect 914 69568 982 69624
rect 1038 69568 1106 69624
rect 1162 69568 1230 69624
rect 1286 69568 1354 69624
rect 1410 69568 1478 69624
rect 1534 69568 1602 69624
rect 1658 69568 1726 69624
rect 1782 69568 1850 69624
rect 1906 69568 2000 69624
rect 0 69500 2000 69568
rect 0 69444 114 69500
rect 170 69444 238 69500
rect 294 69444 362 69500
rect 418 69444 486 69500
rect 542 69444 610 69500
rect 666 69444 734 69500
rect 790 69444 858 69500
rect 914 69444 982 69500
rect 1038 69444 1106 69500
rect 1162 69444 1230 69500
rect 1286 69444 1354 69500
rect 1410 69444 1478 69500
rect 1534 69444 1602 69500
rect 1658 69444 1726 69500
rect 1782 69444 1850 69500
rect 1906 69444 2000 69500
rect 0 69376 2000 69444
rect 0 69320 114 69376
rect 170 69320 238 69376
rect 294 69320 362 69376
rect 418 69320 486 69376
rect 542 69320 610 69376
rect 666 69320 734 69376
rect 790 69320 858 69376
rect 914 69320 982 69376
rect 1038 69320 1106 69376
rect 1162 69320 1230 69376
rect 1286 69320 1354 69376
rect 1410 69320 1478 69376
rect 1534 69320 1602 69376
rect 1658 69320 1726 69376
rect 1782 69320 1850 69376
rect 1906 69320 2000 69376
rect 0 69252 2000 69320
rect 0 69196 114 69252
rect 170 69196 238 69252
rect 294 69196 362 69252
rect 418 69196 486 69252
rect 542 69196 610 69252
rect 666 69196 734 69252
rect 790 69196 858 69252
rect 914 69196 982 69252
rect 1038 69196 1106 69252
rect 1162 69196 1230 69252
rect 1286 69196 1354 69252
rect 1410 69196 1478 69252
rect 1534 69196 1602 69252
rect 1658 69196 1726 69252
rect 1782 69196 1850 69252
rect 1906 69196 2000 69252
rect 0 69128 2000 69196
rect 0 69072 114 69128
rect 170 69072 238 69128
rect 294 69072 362 69128
rect 418 69072 486 69128
rect 542 69072 610 69128
rect 666 69072 734 69128
rect 790 69072 858 69128
rect 914 69072 982 69128
rect 1038 69072 1106 69128
rect 1162 69072 1230 69128
rect 1286 69072 1354 69128
rect 1410 69072 1478 69128
rect 1534 69072 1602 69128
rect 1658 69072 1726 69128
rect 1782 69072 1850 69128
rect 1906 69072 2000 69128
rect 0 69004 2000 69072
rect 0 68948 114 69004
rect 170 68948 238 69004
rect 294 68948 362 69004
rect 418 68948 486 69004
rect 542 68948 610 69004
rect 666 68948 734 69004
rect 790 68948 858 69004
rect 914 68948 982 69004
rect 1038 68948 1106 69004
rect 1162 68948 1230 69004
rect 1286 68948 1354 69004
rect 1410 68948 1478 69004
rect 1534 68948 1602 69004
rect 1658 68948 1726 69004
rect 1782 68948 1850 69004
rect 1906 68948 2000 69004
rect 0 68880 2000 68948
rect 0 68824 114 68880
rect 170 68824 238 68880
rect 294 68824 362 68880
rect 418 68824 486 68880
rect 542 68824 610 68880
rect 666 68824 734 68880
rect 790 68824 858 68880
rect 914 68824 982 68880
rect 1038 68824 1106 68880
rect 1162 68824 1230 68880
rect 1286 68824 1354 68880
rect 1410 68824 1478 68880
rect 1534 68824 1602 68880
rect 1658 68824 1726 68880
rect 1782 68824 1850 68880
rect 1906 68824 2000 68880
rect 0 68756 2000 68824
rect 0 68700 114 68756
rect 170 68700 238 68756
rect 294 68700 362 68756
rect 418 68700 486 68756
rect 542 68700 610 68756
rect 666 68700 734 68756
rect 790 68700 858 68756
rect 914 68700 982 68756
rect 1038 68700 1106 68756
rect 1162 68700 1230 68756
rect 1286 68700 1354 68756
rect 1410 68700 1478 68756
rect 1534 68700 1602 68756
rect 1658 68700 1726 68756
rect 1782 68700 1850 68756
rect 1906 68700 2000 68756
rect 0 68632 2000 68700
rect 0 68576 114 68632
rect 170 68576 238 68632
rect 294 68576 362 68632
rect 418 68576 486 68632
rect 542 68576 610 68632
rect 666 68576 734 68632
rect 790 68576 858 68632
rect 914 68576 982 68632
rect 1038 68576 1106 68632
rect 1162 68576 1230 68632
rect 1286 68576 1354 68632
rect 1410 68576 1478 68632
rect 1534 68576 1602 68632
rect 1658 68576 1726 68632
rect 1782 68576 1850 68632
rect 1906 68576 2000 68632
rect 0 68508 2000 68576
rect 0 68452 114 68508
rect 170 68452 238 68508
rect 294 68452 362 68508
rect 418 68452 486 68508
rect 542 68452 610 68508
rect 666 68452 734 68508
rect 790 68452 858 68508
rect 914 68452 982 68508
rect 1038 68452 1106 68508
rect 1162 68452 1230 68508
rect 1286 68452 1354 68508
rect 1410 68452 1478 68508
rect 1534 68452 1602 68508
rect 1658 68452 1726 68508
rect 1782 68452 1850 68508
rect 1906 68452 2000 68508
rect 0 68400 2000 68452
rect 0 68094 2000 68200
rect 0 68038 114 68094
rect 170 68038 238 68094
rect 294 68038 362 68094
rect 418 68038 486 68094
rect 542 68038 610 68094
rect 666 68038 734 68094
rect 790 68038 858 68094
rect 914 68038 982 68094
rect 1038 68038 1106 68094
rect 1162 68038 1230 68094
rect 1286 68038 1354 68094
rect 1410 68038 1478 68094
rect 1534 68038 1602 68094
rect 1658 68038 1726 68094
rect 1782 68038 1850 68094
rect 1906 68038 2000 68094
rect 0 67970 2000 68038
rect 0 67914 114 67970
rect 170 67914 238 67970
rect 294 67914 362 67970
rect 418 67914 486 67970
rect 542 67914 610 67970
rect 666 67914 734 67970
rect 790 67914 858 67970
rect 914 67914 982 67970
rect 1038 67914 1106 67970
rect 1162 67914 1230 67970
rect 1286 67914 1354 67970
rect 1410 67914 1478 67970
rect 1534 67914 1602 67970
rect 1658 67914 1726 67970
rect 1782 67914 1850 67970
rect 1906 67914 2000 67970
rect 0 67846 2000 67914
rect 0 67790 114 67846
rect 170 67790 238 67846
rect 294 67790 362 67846
rect 418 67790 486 67846
rect 542 67790 610 67846
rect 666 67790 734 67846
rect 790 67790 858 67846
rect 914 67790 982 67846
rect 1038 67790 1106 67846
rect 1162 67790 1230 67846
rect 1286 67790 1354 67846
rect 1410 67790 1478 67846
rect 1534 67790 1602 67846
rect 1658 67790 1726 67846
rect 1782 67790 1850 67846
rect 1906 67790 2000 67846
rect 0 67722 2000 67790
rect 0 67666 114 67722
rect 170 67666 238 67722
rect 294 67666 362 67722
rect 418 67666 486 67722
rect 542 67666 610 67722
rect 666 67666 734 67722
rect 790 67666 858 67722
rect 914 67666 982 67722
rect 1038 67666 1106 67722
rect 1162 67666 1230 67722
rect 1286 67666 1354 67722
rect 1410 67666 1478 67722
rect 1534 67666 1602 67722
rect 1658 67666 1726 67722
rect 1782 67666 1850 67722
rect 1906 67666 2000 67722
rect 0 67598 2000 67666
rect 0 67542 114 67598
rect 170 67542 238 67598
rect 294 67542 362 67598
rect 418 67542 486 67598
rect 542 67542 610 67598
rect 666 67542 734 67598
rect 790 67542 858 67598
rect 914 67542 982 67598
rect 1038 67542 1106 67598
rect 1162 67542 1230 67598
rect 1286 67542 1354 67598
rect 1410 67542 1478 67598
rect 1534 67542 1602 67598
rect 1658 67542 1726 67598
rect 1782 67542 1850 67598
rect 1906 67542 2000 67598
rect 0 67474 2000 67542
rect 0 67418 114 67474
rect 170 67418 238 67474
rect 294 67418 362 67474
rect 418 67418 486 67474
rect 542 67418 610 67474
rect 666 67418 734 67474
rect 790 67418 858 67474
rect 914 67418 982 67474
rect 1038 67418 1106 67474
rect 1162 67418 1230 67474
rect 1286 67418 1354 67474
rect 1410 67418 1478 67474
rect 1534 67418 1602 67474
rect 1658 67418 1726 67474
rect 1782 67418 1850 67474
rect 1906 67418 2000 67474
rect 0 67350 2000 67418
rect 0 67294 114 67350
rect 170 67294 238 67350
rect 294 67294 362 67350
rect 418 67294 486 67350
rect 542 67294 610 67350
rect 666 67294 734 67350
rect 790 67294 858 67350
rect 914 67294 982 67350
rect 1038 67294 1106 67350
rect 1162 67294 1230 67350
rect 1286 67294 1354 67350
rect 1410 67294 1478 67350
rect 1534 67294 1602 67350
rect 1658 67294 1726 67350
rect 1782 67294 1850 67350
rect 1906 67294 2000 67350
rect 0 67226 2000 67294
rect 0 67170 114 67226
rect 170 67170 238 67226
rect 294 67170 362 67226
rect 418 67170 486 67226
rect 542 67170 610 67226
rect 666 67170 734 67226
rect 790 67170 858 67226
rect 914 67170 982 67226
rect 1038 67170 1106 67226
rect 1162 67170 1230 67226
rect 1286 67170 1354 67226
rect 1410 67170 1478 67226
rect 1534 67170 1602 67226
rect 1658 67170 1726 67226
rect 1782 67170 1850 67226
rect 1906 67170 2000 67226
rect 0 67102 2000 67170
rect 0 67046 114 67102
rect 170 67046 238 67102
rect 294 67046 362 67102
rect 418 67046 486 67102
rect 542 67046 610 67102
rect 666 67046 734 67102
rect 790 67046 858 67102
rect 914 67046 982 67102
rect 1038 67046 1106 67102
rect 1162 67046 1230 67102
rect 1286 67046 1354 67102
rect 1410 67046 1478 67102
rect 1534 67046 1602 67102
rect 1658 67046 1726 67102
rect 1782 67046 1850 67102
rect 1906 67046 2000 67102
rect 0 66978 2000 67046
rect 0 66922 114 66978
rect 170 66922 238 66978
rect 294 66922 362 66978
rect 418 66922 486 66978
rect 542 66922 610 66978
rect 666 66922 734 66978
rect 790 66922 858 66978
rect 914 66922 982 66978
rect 1038 66922 1106 66978
rect 1162 66922 1230 66978
rect 1286 66922 1354 66978
rect 1410 66922 1478 66978
rect 1534 66922 1602 66978
rect 1658 66922 1726 66978
rect 1782 66922 1850 66978
rect 1906 66922 2000 66978
rect 0 66800 2000 66922
rect 0 66484 2000 66600
rect 0 66428 114 66484
rect 170 66428 238 66484
rect 294 66428 362 66484
rect 418 66428 486 66484
rect 542 66428 610 66484
rect 666 66428 734 66484
rect 790 66428 858 66484
rect 914 66428 982 66484
rect 1038 66428 1106 66484
rect 1162 66428 1230 66484
rect 1286 66428 1354 66484
rect 1410 66428 1478 66484
rect 1534 66428 1602 66484
rect 1658 66428 1726 66484
rect 1782 66428 1850 66484
rect 1906 66428 2000 66484
rect 0 66360 2000 66428
rect 0 66304 114 66360
rect 170 66304 238 66360
rect 294 66304 362 66360
rect 418 66304 486 66360
rect 542 66304 610 66360
rect 666 66304 734 66360
rect 790 66304 858 66360
rect 914 66304 982 66360
rect 1038 66304 1106 66360
rect 1162 66304 1230 66360
rect 1286 66304 1354 66360
rect 1410 66304 1478 66360
rect 1534 66304 1602 66360
rect 1658 66304 1726 66360
rect 1782 66304 1850 66360
rect 1906 66304 2000 66360
rect 0 66236 2000 66304
rect 0 66180 114 66236
rect 170 66180 238 66236
rect 294 66180 362 66236
rect 418 66180 486 66236
rect 542 66180 610 66236
rect 666 66180 734 66236
rect 790 66180 858 66236
rect 914 66180 982 66236
rect 1038 66180 1106 66236
rect 1162 66180 1230 66236
rect 1286 66180 1354 66236
rect 1410 66180 1478 66236
rect 1534 66180 1602 66236
rect 1658 66180 1726 66236
rect 1782 66180 1850 66236
rect 1906 66180 2000 66236
rect 0 66112 2000 66180
rect 0 66056 114 66112
rect 170 66056 238 66112
rect 294 66056 362 66112
rect 418 66056 486 66112
rect 542 66056 610 66112
rect 666 66056 734 66112
rect 790 66056 858 66112
rect 914 66056 982 66112
rect 1038 66056 1106 66112
rect 1162 66056 1230 66112
rect 1286 66056 1354 66112
rect 1410 66056 1478 66112
rect 1534 66056 1602 66112
rect 1658 66056 1726 66112
rect 1782 66056 1850 66112
rect 1906 66056 2000 66112
rect 0 65988 2000 66056
rect 0 65932 114 65988
rect 170 65932 238 65988
rect 294 65932 362 65988
rect 418 65932 486 65988
rect 542 65932 610 65988
rect 666 65932 734 65988
rect 790 65932 858 65988
rect 914 65932 982 65988
rect 1038 65932 1106 65988
rect 1162 65932 1230 65988
rect 1286 65932 1354 65988
rect 1410 65932 1478 65988
rect 1534 65932 1602 65988
rect 1658 65932 1726 65988
rect 1782 65932 1850 65988
rect 1906 65932 2000 65988
rect 0 65864 2000 65932
rect 0 65808 114 65864
rect 170 65808 238 65864
rect 294 65808 362 65864
rect 418 65808 486 65864
rect 542 65808 610 65864
rect 666 65808 734 65864
rect 790 65808 858 65864
rect 914 65808 982 65864
rect 1038 65808 1106 65864
rect 1162 65808 1230 65864
rect 1286 65808 1354 65864
rect 1410 65808 1478 65864
rect 1534 65808 1602 65864
rect 1658 65808 1726 65864
rect 1782 65808 1850 65864
rect 1906 65808 2000 65864
rect 0 65740 2000 65808
rect 0 65684 114 65740
rect 170 65684 238 65740
rect 294 65684 362 65740
rect 418 65684 486 65740
rect 542 65684 610 65740
rect 666 65684 734 65740
rect 790 65684 858 65740
rect 914 65684 982 65740
rect 1038 65684 1106 65740
rect 1162 65684 1230 65740
rect 1286 65684 1354 65740
rect 1410 65684 1478 65740
rect 1534 65684 1602 65740
rect 1658 65684 1726 65740
rect 1782 65684 1850 65740
rect 1906 65684 2000 65740
rect 0 65616 2000 65684
rect 0 65560 114 65616
rect 170 65560 238 65616
rect 294 65560 362 65616
rect 418 65560 486 65616
rect 542 65560 610 65616
rect 666 65560 734 65616
rect 790 65560 858 65616
rect 914 65560 982 65616
rect 1038 65560 1106 65616
rect 1162 65560 1230 65616
rect 1286 65560 1354 65616
rect 1410 65560 1478 65616
rect 1534 65560 1602 65616
rect 1658 65560 1726 65616
rect 1782 65560 1850 65616
rect 1906 65560 2000 65616
rect 0 65492 2000 65560
rect 0 65436 114 65492
rect 170 65436 238 65492
rect 294 65436 362 65492
rect 418 65436 486 65492
rect 542 65436 610 65492
rect 666 65436 734 65492
rect 790 65436 858 65492
rect 914 65436 982 65492
rect 1038 65436 1106 65492
rect 1162 65436 1230 65492
rect 1286 65436 1354 65492
rect 1410 65436 1478 65492
rect 1534 65436 1602 65492
rect 1658 65436 1726 65492
rect 1782 65436 1850 65492
rect 1906 65436 2000 65492
rect 0 65368 2000 65436
rect 0 65312 114 65368
rect 170 65312 238 65368
rect 294 65312 362 65368
rect 418 65312 486 65368
rect 542 65312 610 65368
rect 666 65312 734 65368
rect 790 65312 858 65368
rect 914 65312 982 65368
rect 1038 65312 1106 65368
rect 1162 65312 1230 65368
rect 1286 65312 1354 65368
rect 1410 65312 1478 65368
rect 1534 65312 1602 65368
rect 1658 65312 1726 65368
rect 1782 65312 1850 65368
rect 1906 65312 2000 65368
rect 0 65200 2000 65312
rect 0 64886 2000 65000
rect 0 64830 114 64886
rect 170 64830 238 64886
rect 294 64830 362 64886
rect 418 64830 486 64886
rect 542 64830 610 64886
rect 666 64830 734 64886
rect 790 64830 858 64886
rect 914 64830 982 64886
rect 1038 64830 1106 64886
rect 1162 64830 1230 64886
rect 1286 64830 1354 64886
rect 1410 64830 1478 64886
rect 1534 64830 1602 64886
rect 1658 64830 1726 64886
rect 1782 64830 1850 64886
rect 1906 64830 2000 64886
rect 0 64762 2000 64830
rect 0 64706 114 64762
rect 170 64706 238 64762
rect 294 64706 362 64762
rect 418 64706 486 64762
rect 542 64706 610 64762
rect 666 64706 734 64762
rect 790 64706 858 64762
rect 914 64706 982 64762
rect 1038 64706 1106 64762
rect 1162 64706 1230 64762
rect 1286 64706 1354 64762
rect 1410 64706 1478 64762
rect 1534 64706 1602 64762
rect 1658 64706 1726 64762
rect 1782 64706 1850 64762
rect 1906 64706 2000 64762
rect 0 64638 2000 64706
rect 0 64582 114 64638
rect 170 64582 238 64638
rect 294 64582 362 64638
rect 418 64582 486 64638
rect 542 64582 610 64638
rect 666 64582 734 64638
rect 790 64582 858 64638
rect 914 64582 982 64638
rect 1038 64582 1106 64638
rect 1162 64582 1230 64638
rect 1286 64582 1354 64638
rect 1410 64582 1478 64638
rect 1534 64582 1602 64638
rect 1658 64582 1726 64638
rect 1782 64582 1850 64638
rect 1906 64582 2000 64638
rect 0 64514 2000 64582
rect 0 64458 114 64514
rect 170 64458 238 64514
rect 294 64458 362 64514
rect 418 64458 486 64514
rect 542 64458 610 64514
rect 666 64458 734 64514
rect 790 64458 858 64514
rect 914 64458 982 64514
rect 1038 64458 1106 64514
rect 1162 64458 1230 64514
rect 1286 64458 1354 64514
rect 1410 64458 1478 64514
rect 1534 64458 1602 64514
rect 1658 64458 1726 64514
rect 1782 64458 1850 64514
rect 1906 64458 2000 64514
rect 0 64390 2000 64458
rect 0 64334 114 64390
rect 170 64334 238 64390
rect 294 64334 362 64390
rect 418 64334 486 64390
rect 542 64334 610 64390
rect 666 64334 734 64390
rect 790 64334 858 64390
rect 914 64334 982 64390
rect 1038 64334 1106 64390
rect 1162 64334 1230 64390
rect 1286 64334 1354 64390
rect 1410 64334 1478 64390
rect 1534 64334 1602 64390
rect 1658 64334 1726 64390
rect 1782 64334 1850 64390
rect 1906 64334 2000 64390
rect 0 64266 2000 64334
rect 0 64210 114 64266
rect 170 64210 238 64266
rect 294 64210 362 64266
rect 418 64210 486 64266
rect 542 64210 610 64266
rect 666 64210 734 64266
rect 790 64210 858 64266
rect 914 64210 982 64266
rect 1038 64210 1106 64266
rect 1162 64210 1230 64266
rect 1286 64210 1354 64266
rect 1410 64210 1478 64266
rect 1534 64210 1602 64266
rect 1658 64210 1726 64266
rect 1782 64210 1850 64266
rect 1906 64210 2000 64266
rect 0 64142 2000 64210
rect 0 64086 114 64142
rect 170 64086 238 64142
rect 294 64086 362 64142
rect 418 64086 486 64142
rect 542 64086 610 64142
rect 666 64086 734 64142
rect 790 64086 858 64142
rect 914 64086 982 64142
rect 1038 64086 1106 64142
rect 1162 64086 1230 64142
rect 1286 64086 1354 64142
rect 1410 64086 1478 64142
rect 1534 64086 1602 64142
rect 1658 64086 1726 64142
rect 1782 64086 1850 64142
rect 1906 64086 2000 64142
rect 0 64018 2000 64086
rect 0 63962 114 64018
rect 170 63962 238 64018
rect 294 63962 362 64018
rect 418 63962 486 64018
rect 542 63962 610 64018
rect 666 63962 734 64018
rect 790 63962 858 64018
rect 914 63962 982 64018
rect 1038 63962 1106 64018
rect 1162 63962 1230 64018
rect 1286 63962 1354 64018
rect 1410 63962 1478 64018
rect 1534 63962 1602 64018
rect 1658 63962 1726 64018
rect 1782 63962 1850 64018
rect 1906 63962 2000 64018
rect 0 63894 2000 63962
rect 0 63838 114 63894
rect 170 63838 238 63894
rect 294 63838 362 63894
rect 418 63838 486 63894
rect 542 63838 610 63894
rect 666 63838 734 63894
rect 790 63838 858 63894
rect 914 63838 982 63894
rect 1038 63838 1106 63894
rect 1162 63838 1230 63894
rect 1286 63838 1354 63894
rect 1410 63838 1478 63894
rect 1534 63838 1602 63894
rect 1658 63838 1726 63894
rect 1782 63838 1850 63894
rect 1906 63838 2000 63894
rect 0 63770 2000 63838
rect 0 63714 114 63770
rect 170 63714 238 63770
rect 294 63714 362 63770
rect 418 63714 486 63770
rect 542 63714 610 63770
rect 666 63714 734 63770
rect 790 63714 858 63770
rect 914 63714 982 63770
rect 1038 63714 1106 63770
rect 1162 63714 1230 63770
rect 1286 63714 1354 63770
rect 1410 63714 1478 63770
rect 1534 63714 1602 63770
rect 1658 63714 1726 63770
rect 1782 63714 1850 63770
rect 1906 63714 2000 63770
rect 0 63600 2000 63714
rect 0 63295 2000 63400
rect 0 63239 114 63295
rect 170 63239 238 63295
rect 294 63239 362 63295
rect 418 63239 486 63295
rect 542 63239 610 63295
rect 666 63239 734 63295
rect 790 63239 858 63295
rect 914 63239 982 63295
rect 1038 63239 1106 63295
rect 1162 63239 1230 63295
rect 1286 63239 1354 63295
rect 1410 63239 1478 63295
rect 1534 63239 1602 63295
rect 1658 63239 1726 63295
rect 1782 63239 1850 63295
rect 1906 63239 2000 63295
rect 0 63171 2000 63239
rect 0 63115 114 63171
rect 170 63115 238 63171
rect 294 63115 362 63171
rect 418 63115 486 63171
rect 542 63115 610 63171
rect 666 63115 734 63171
rect 790 63115 858 63171
rect 914 63115 982 63171
rect 1038 63115 1106 63171
rect 1162 63115 1230 63171
rect 1286 63115 1354 63171
rect 1410 63115 1478 63171
rect 1534 63115 1602 63171
rect 1658 63115 1726 63171
rect 1782 63115 1850 63171
rect 1906 63115 2000 63171
rect 0 63047 2000 63115
rect 0 62991 114 63047
rect 170 62991 238 63047
rect 294 62991 362 63047
rect 418 62991 486 63047
rect 542 62991 610 63047
rect 666 62991 734 63047
rect 790 62991 858 63047
rect 914 62991 982 63047
rect 1038 62991 1106 63047
rect 1162 62991 1230 63047
rect 1286 62991 1354 63047
rect 1410 62991 1478 63047
rect 1534 62991 1602 63047
rect 1658 62991 1726 63047
rect 1782 62991 1850 63047
rect 1906 62991 2000 63047
rect 0 62923 2000 62991
rect 0 62867 114 62923
rect 170 62867 238 62923
rect 294 62867 362 62923
rect 418 62867 486 62923
rect 542 62867 610 62923
rect 666 62867 734 62923
rect 790 62867 858 62923
rect 914 62867 982 62923
rect 1038 62867 1106 62923
rect 1162 62867 1230 62923
rect 1286 62867 1354 62923
rect 1410 62867 1478 62923
rect 1534 62867 1602 62923
rect 1658 62867 1726 62923
rect 1782 62867 1850 62923
rect 1906 62867 2000 62923
rect 0 62799 2000 62867
rect 0 62743 114 62799
rect 170 62743 238 62799
rect 294 62743 362 62799
rect 418 62743 486 62799
rect 542 62743 610 62799
rect 666 62743 734 62799
rect 790 62743 858 62799
rect 914 62743 982 62799
rect 1038 62743 1106 62799
rect 1162 62743 1230 62799
rect 1286 62743 1354 62799
rect 1410 62743 1478 62799
rect 1534 62743 1602 62799
rect 1658 62743 1726 62799
rect 1782 62743 1850 62799
rect 1906 62743 2000 62799
rect 0 62675 2000 62743
rect 0 62619 114 62675
rect 170 62619 238 62675
rect 294 62619 362 62675
rect 418 62619 486 62675
rect 542 62619 610 62675
rect 666 62619 734 62675
rect 790 62619 858 62675
rect 914 62619 982 62675
rect 1038 62619 1106 62675
rect 1162 62619 1230 62675
rect 1286 62619 1354 62675
rect 1410 62619 1478 62675
rect 1534 62619 1602 62675
rect 1658 62619 1726 62675
rect 1782 62619 1850 62675
rect 1906 62619 2000 62675
rect 0 62551 2000 62619
rect 0 62495 114 62551
rect 170 62495 238 62551
rect 294 62495 362 62551
rect 418 62495 486 62551
rect 542 62495 610 62551
rect 666 62495 734 62551
rect 790 62495 858 62551
rect 914 62495 982 62551
rect 1038 62495 1106 62551
rect 1162 62495 1230 62551
rect 1286 62495 1354 62551
rect 1410 62495 1478 62551
rect 1534 62495 1602 62551
rect 1658 62495 1726 62551
rect 1782 62495 1850 62551
rect 1906 62495 2000 62551
rect 0 62427 2000 62495
rect 0 62371 114 62427
rect 170 62371 238 62427
rect 294 62371 362 62427
rect 418 62371 486 62427
rect 542 62371 610 62427
rect 666 62371 734 62427
rect 790 62371 858 62427
rect 914 62371 982 62427
rect 1038 62371 1106 62427
rect 1162 62371 1230 62427
rect 1286 62371 1354 62427
rect 1410 62371 1478 62427
rect 1534 62371 1602 62427
rect 1658 62371 1726 62427
rect 1782 62371 1850 62427
rect 1906 62371 2000 62427
rect 0 62303 2000 62371
rect 0 62247 114 62303
rect 170 62247 238 62303
rect 294 62247 362 62303
rect 418 62247 486 62303
rect 542 62247 610 62303
rect 666 62247 734 62303
rect 790 62247 858 62303
rect 914 62247 982 62303
rect 1038 62247 1106 62303
rect 1162 62247 1230 62303
rect 1286 62247 1354 62303
rect 1410 62247 1478 62303
rect 1534 62247 1602 62303
rect 1658 62247 1726 62303
rect 1782 62247 1850 62303
rect 1906 62247 2000 62303
rect 0 62179 2000 62247
rect 0 62123 114 62179
rect 170 62123 238 62179
rect 294 62123 362 62179
rect 418 62123 486 62179
rect 542 62123 610 62179
rect 666 62123 734 62179
rect 790 62123 858 62179
rect 914 62123 982 62179
rect 1038 62123 1106 62179
rect 1162 62123 1230 62179
rect 1286 62123 1354 62179
rect 1410 62123 1478 62179
rect 1534 62123 1602 62179
rect 1658 62123 1726 62179
rect 1782 62123 1850 62179
rect 1906 62123 2000 62179
rect 0 62000 2000 62123
rect 0 61695 2000 61800
rect 0 61639 114 61695
rect 170 61639 238 61695
rect 294 61639 362 61695
rect 418 61639 486 61695
rect 542 61639 610 61695
rect 666 61639 734 61695
rect 790 61639 858 61695
rect 914 61639 982 61695
rect 1038 61639 1106 61695
rect 1162 61639 1230 61695
rect 1286 61639 1354 61695
rect 1410 61639 1478 61695
rect 1534 61639 1602 61695
rect 1658 61639 1726 61695
rect 1782 61639 1850 61695
rect 1906 61639 2000 61695
rect 0 61571 2000 61639
rect 0 61515 114 61571
rect 170 61515 238 61571
rect 294 61515 362 61571
rect 418 61515 486 61571
rect 542 61515 610 61571
rect 666 61515 734 61571
rect 790 61515 858 61571
rect 914 61515 982 61571
rect 1038 61515 1106 61571
rect 1162 61515 1230 61571
rect 1286 61515 1354 61571
rect 1410 61515 1478 61571
rect 1534 61515 1602 61571
rect 1658 61515 1726 61571
rect 1782 61515 1850 61571
rect 1906 61515 2000 61571
rect 0 61447 2000 61515
rect 0 61391 114 61447
rect 170 61391 238 61447
rect 294 61391 362 61447
rect 418 61391 486 61447
rect 542 61391 610 61447
rect 666 61391 734 61447
rect 790 61391 858 61447
rect 914 61391 982 61447
rect 1038 61391 1106 61447
rect 1162 61391 1230 61447
rect 1286 61391 1354 61447
rect 1410 61391 1478 61447
rect 1534 61391 1602 61447
rect 1658 61391 1726 61447
rect 1782 61391 1850 61447
rect 1906 61391 2000 61447
rect 0 61323 2000 61391
rect 0 61267 114 61323
rect 170 61267 238 61323
rect 294 61267 362 61323
rect 418 61267 486 61323
rect 542 61267 610 61323
rect 666 61267 734 61323
rect 790 61267 858 61323
rect 914 61267 982 61323
rect 1038 61267 1106 61323
rect 1162 61267 1230 61323
rect 1286 61267 1354 61323
rect 1410 61267 1478 61323
rect 1534 61267 1602 61323
rect 1658 61267 1726 61323
rect 1782 61267 1850 61323
rect 1906 61267 2000 61323
rect 0 61199 2000 61267
rect 0 61143 114 61199
rect 170 61143 238 61199
rect 294 61143 362 61199
rect 418 61143 486 61199
rect 542 61143 610 61199
rect 666 61143 734 61199
rect 790 61143 858 61199
rect 914 61143 982 61199
rect 1038 61143 1106 61199
rect 1162 61143 1230 61199
rect 1286 61143 1354 61199
rect 1410 61143 1478 61199
rect 1534 61143 1602 61199
rect 1658 61143 1726 61199
rect 1782 61143 1850 61199
rect 1906 61143 2000 61199
rect 0 61075 2000 61143
rect 0 61019 114 61075
rect 170 61019 238 61075
rect 294 61019 362 61075
rect 418 61019 486 61075
rect 542 61019 610 61075
rect 666 61019 734 61075
rect 790 61019 858 61075
rect 914 61019 982 61075
rect 1038 61019 1106 61075
rect 1162 61019 1230 61075
rect 1286 61019 1354 61075
rect 1410 61019 1478 61075
rect 1534 61019 1602 61075
rect 1658 61019 1726 61075
rect 1782 61019 1850 61075
rect 1906 61019 2000 61075
rect 0 60951 2000 61019
rect 0 60895 114 60951
rect 170 60895 238 60951
rect 294 60895 362 60951
rect 418 60895 486 60951
rect 542 60895 610 60951
rect 666 60895 734 60951
rect 790 60895 858 60951
rect 914 60895 982 60951
rect 1038 60895 1106 60951
rect 1162 60895 1230 60951
rect 1286 60895 1354 60951
rect 1410 60895 1478 60951
rect 1534 60895 1602 60951
rect 1658 60895 1726 60951
rect 1782 60895 1850 60951
rect 1906 60895 2000 60951
rect 0 60827 2000 60895
rect 0 60771 114 60827
rect 170 60771 238 60827
rect 294 60771 362 60827
rect 418 60771 486 60827
rect 542 60771 610 60827
rect 666 60771 734 60827
rect 790 60771 858 60827
rect 914 60771 982 60827
rect 1038 60771 1106 60827
rect 1162 60771 1230 60827
rect 1286 60771 1354 60827
rect 1410 60771 1478 60827
rect 1534 60771 1602 60827
rect 1658 60771 1726 60827
rect 1782 60771 1850 60827
rect 1906 60771 2000 60827
rect 0 60703 2000 60771
rect 0 60647 114 60703
rect 170 60647 238 60703
rect 294 60647 362 60703
rect 418 60647 486 60703
rect 542 60647 610 60703
rect 666 60647 734 60703
rect 790 60647 858 60703
rect 914 60647 982 60703
rect 1038 60647 1106 60703
rect 1162 60647 1230 60703
rect 1286 60647 1354 60703
rect 1410 60647 1478 60703
rect 1534 60647 1602 60703
rect 1658 60647 1726 60703
rect 1782 60647 1850 60703
rect 1906 60647 2000 60703
rect 0 60579 2000 60647
rect 0 60523 114 60579
rect 170 60523 238 60579
rect 294 60523 362 60579
rect 418 60523 486 60579
rect 542 60523 610 60579
rect 666 60523 734 60579
rect 790 60523 858 60579
rect 914 60523 982 60579
rect 1038 60523 1106 60579
rect 1162 60523 1230 60579
rect 1286 60523 1354 60579
rect 1410 60523 1478 60579
rect 1534 60523 1602 60579
rect 1658 60523 1726 60579
rect 1782 60523 1850 60579
rect 1906 60523 2000 60579
rect 0 60400 2000 60523
rect 0 60090 2000 60200
rect 0 60034 114 60090
rect 170 60034 238 60090
rect 294 60034 362 60090
rect 418 60034 486 60090
rect 542 60034 610 60090
rect 666 60034 734 60090
rect 790 60034 858 60090
rect 914 60034 982 60090
rect 1038 60034 1106 60090
rect 1162 60034 1230 60090
rect 1286 60034 1354 60090
rect 1410 60034 1478 60090
rect 1534 60034 1602 60090
rect 1658 60034 1726 60090
rect 1782 60034 1850 60090
rect 1906 60034 2000 60090
rect 0 59966 2000 60034
rect 0 59910 114 59966
rect 170 59910 238 59966
rect 294 59910 362 59966
rect 418 59910 486 59966
rect 542 59910 610 59966
rect 666 59910 734 59966
rect 790 59910 858 59966
rect 914 59910 982 59966
rect 1038 59910 1106 59966
rect 1162 59910 1230 59966
rect 1286 59910 1354 59966
rect 1410 59910 1478 59966
rect 1534 59910 1602 59966
rect 1658 59910 1726 59966
rect 1782 59910 1850 59966
rect 1906 59910 2000 59966
rect 0 59842 2000 59910
rect 0 59786 114 59842
rect 170 59786 238 59842
rect 294 59786 362 59842
rect 418 59786 486 59842
rect 542 59786 610 59842
rect 666 59786 734 59842
rect 790 59786 858 59842
rect 914 59786 982 59842
rect 1038 59786 1106 59842
rect 1162 59786 1230 59842
rect 1286 59786 1354 59842
rect 1410 59786 1478 59842
rect 1534 59786 1602 59842
rect 1658 59786 1726 59842
rect 1782 59786 1850 59842
rect 1906 59786 2000 59842
rect 0 59718 2000 59786
rect 0 59662 114 59718
rect 170 59662 238 59718
rect 294 59662 362 59718
rect 418 59662 486 59718
rect 542 59662 610 59718
rect 666 59662 734 59718
rect 790 59662 858 59718
rect 914 59662 982 59718
rect 1038 59662 1106 59718
rect 1162 59662 1230 59718
rect 1286 59662 1354 59718
rect 1410 59662 1478 59718
rect 1534 59662 1602 59718
rect 1658 59662 1726 59718
rect 1782 59662 1850 59718
rect 1906 59662 2000 59718
rect 0 59594 2000 59662
rect 0 59538 114 59594
rect 170 59538 238 59594
rect 294 59538 362 59594
rect 418 59538 486 59594
rect 542 59538 610 59594
rect 666 59538 734 59594
rect 790 59538 858 59594
rect 914 59538 982 59594
rect 1038 59538 1106 59594
rect 1162 59538 1230 59594
rect 1286 59538 1354 59594
rect 1410 59538 1478 59594
rect 1534 59538 1602 59594
rect 1658 59538 1726 59594
rect 1782 59538 1850 59594
rect 1906 59538 2000 59594
rect 0 59470 2000 59538
rect 0 59414 114 59470
rect 170 59414 238 59470
rect 294 59414 362 59470
rect 418 59414 486 59470
rect 542 59414 610 59470
rect 666 59414 734 59470
rect 790 59414 858 59470
rect 914 59414 982 59470
rect 1038 59414 1106 59470
rect 1162 59414 1230 59470
rect 1286 59414 1354 59470
rect 1410 59414 1478 59470
rect 1534 59414 1602 59470
rect 1658 59414 1726 59470
rect 1782 59414 1850 59470
rect 1906 59414 2000 59470
rect 0 59346 2000 59414
rect 0 59290 114 59346
rect 170 59290 238 59346
rect 294 59290 362 59346
rect 418 59290 486 59346
rect 542 59290 610 59346
rect 666 59290 734 59346
rect 790 59290 858 59346
rect 914 59290 982 59346
rect 1038 59290 1106 59346
rect 1162 59290 1230 59346
rect 1286 59290 1354 59346
rect 1410 59290 1478 59346
rect 1534 59290 1602 59346
rect 1658 59290 1726 59346
rect 1782 59290 1850 59346
rect 1906 59290 2000 59346
rect 0 59222 2000 59290
rect 0 59166 114 59222
rect 170 59166 238 59222
rect 294 59166 362 59222
rect 418 59166 486 59222
rect 542 59166 610 59222
rect 666 59166 734 59222
rect 790 59166 858 59222
rect 914 59166 982 59222
rect 1038 59166 1106 59222
rect 1162 59166 1230 59222
rect 1286 59166 1354 59222
rect 1410 59166 1478 59222
rect 1534 59166 1602 59222
rect 1658 59166 1726 59222
rect 1782 59166 1850 59222
rect 1906 59166 2000 59222
rect 0 59098 2000 59166
rect 0 59042 114 59098
rect 170 59042 238 59098
rect 294 59042 362 59098
rect 418 59042 486 59098
rect 542 59042 610 59098
rect 666 59042 734 59098
rect 790 59042 858 59098
rect 914 59042 982 59098
rect 1038 59042 1106 59098
rect 1162 59042 1230 59098
rect 1286 59042 1354 59098
rect 1410 59042 1478 59098
rect 1534 59042 1602 59098
rect 1658 59042 1726 59098
rect 1782 59042 1850 59098
rect 1906 59042 2000 59098
rect 0 58974 2000 59042
rect 0 58918 114 58974
rect 170 58918 238 58974
rect 294 58918 362 58974
rect 418 58918 486 58974
rect 542 58918 610 58974
rect 666 58918 734 58974
rect 790 58918 858 58974
rect 914 58918 982 58974
rect 1038 58918 1106 58974
rect 1162 58918 1230 58974
rect 1286 58918 1354 58974
rect 1410 58918 1478 58974
rect 1534 58918 1602 58974
rect 1658 58918 1726 58974
rect 1782 58918 1850 58974
rect 1906 58918 2000 58974
rect 0 58800 2000 58918
rect 0 58485 2000 58600
rect 0 58429 114 58485
rect 170 58429 238 58485
rect 294 58429 362 58485
rect 418 58429 486 58485
rect 542 58429 610 58485
rect 666 58429 734 58485
rect 790 58429 858 58485
rect 914 58429 982 58485
rect 1038 58429 1106 58485
rect 1162 58429 1230 58485
rect 1286 58429 1354 58485
rect 1410 58429 1478 58485
rect 1534 58429 1602 58485
rect 1658 58429 1726 58485
rect 1782 58429 1850 58485
rect 1906 58429 2000 58485
rect 0 58361 2000 58429
rect 0 58305 114 58361
rect 170 58305 238 58361
rect 294 58305 362 58361
rect 418 58305 486 58361
rect 542 58305 610 58361
rect 666 58305 734 58361
rect 790 58305 858 58361
rect 914 58305 982 58361
rect 1038 58305 1106 58361
rect 1162 58305 1230 58361
rect 1286 58305 1354 58361
rect 1410 58305 1478 58361
rect 1534 58305 1602 58361
rect 1658 58305 1726 58361
rect 1782 58305 1850 58361
rect 1906 58305 2000 58361
rect 0 58237 2000 58305
rect 0 58181 114 58237
rect 170 58181 238 58237
rect 294 58181 362 58237
rect 418 58181 486 58237
rect 542 58181 610 58237
rect 666 58181 734 58237
rect 790 58181 858 58237
rect 914 58181 982 58237
rect 1038 58181 1106 58237
rect 1162 58181 1230 58237
rect 1286 58181 1354 58237
rect 1410 58181 1478 58237
rect 1534 58181 1602 58237
rect 1658 58181 1726 58237
rect 1782 58181 1850 58237
rect 1906 58181 2000 58237
rect 0 58113 2000 58181
rect 0 58057 114 58113
rect 170 58057 238 58113
rect 294 58057 362 58113
rect 418 58057 486 58113
rect 542 58057 610 58113
rect 666 58057 734 58113
rect 790 58057 858 58113
rect 914 58057 982 58113
rect 1038 58057 1106 58113
rect 1162 58057 1230 58113
rect 1286 58057 1354 58113
rect 1410 58057 1478 58113
rect 1534 58057 1602 58113
rect 1658 58057 1726 58113
rect 1782 58057 1850 58113
rect 1906 58057 2000 58113
rect 0 57989 2000 58057
rect 0 57933 114 57989
rect 170 57933 238 57989
rect 294 57933 362 57989
rect 418 57933 486 57989
rect 542 57933 610 57989
rect 666 57933 734 57989
rect 790 57933 858 57989
rect 914 57933 982 57989
rect 1038 57933 1106 57989
rect 1162 57933 1230 57989
rect 1286 57933 1354 57989
rect 1410 57933 1478 57989
rect 1534 57933 1602 57989
rect 1658 57933 1726 57989
rect 1782 57933 1850 57989
rect 1906 57933 2000 57989
rect 0 57865 2000 57933
rect 0 57809 114 57865
rect 170 57809 238 57865
rect 294 57809 362 57865
rect 418 57809 486 57865
rect 542 57809 610 57865
rect 666 57809 734 57865
rect 790 57809 858 57865
rect 914 57809 982 57865
rect 1038 57809 1106 57865
rect 1162 57809 1230 57865
rect 1286 57809 1354 57865
rect 1410 57809 1478 57865
rect 1534 57809 1602 57865
rect 1658 57809 1726 57865
rect 1782 57809 1850 57865
rect 1906 57809 2000 57865
rect 0 57741 2000 57809
rect 0 57685 114 57741
rect 170 57685 238 57741
rect 294 57685 362 57741
rect 418 57685 486 57741
rect 542 57685 610 57741
rect 666 57685 734 57741
rect 790 57685 858 57741
rect 914 57685 982 57741
rect 1038 57685 1106 57741
rect 1162 57685 1230 57741
rect 1286 57685 1354 57741
rect 1410 57685 1478 57741
rect 1534 57685 1602 57741
rect 1658 57685 1726 57741
rect 1782 57685 1850 57741
rect 1906 57685 2000 57741
rect 0 57617 2000 57685
rect 0 57561 114 57617
rect 170 57561 238 57617
rect 294 57561 362 57617
rect 418 57561 486 57617
rect 542 57561 610 57617
rect 666 57561 734 57617
rect 790 57561 858 57617
rect 914 57561 982 57617
rect 1038 57561 1106 57617
rect 1162 57561 1230 57617
rect 1286 57561 1354 57617
rect 1410 57561 1478 57617
rect 1534 57561 1602 57617
rect 1658 57561 1726 57617
rect 1782 57561 1850 57617
rect 1906 57561 2000 57617
rect 0 57493 2000 57561
rect 0 57437 114 57493
rect 170 57437 238 57493
rect 294 57437 362 57493
rect 418 57437 486 57493
rect 542 57437 610 57493
rect 666 57437 734 57493
rect 790 57437 858 57493
rect 914 57437 982 57493
rect 1038 57437 1106 57493
rect 1162 57437 1230 57493
rect 1286 57437 1354 57493
rect 1410 57437 1478 57493
rect 1534 57437 1602 57493
rect 1658 57437 1726 57493
rect 1782 57437 1850 57493
rect 1906 57437 2000 57493
rect 0 57369 2000 57437
rect 0 57313 114 57369
rect 170 57313 238 57369
rect 294 57313 362 57369
rect 418 57313 486 57369
rect 542 57313 610 57369
rect 666 57313 734 57369
rect 790 57313 858 57369
rect 914 57313 982 57369
rect 1038 57313 1106 57369
rect 1162 57313 1230 57369
rect 1286 57313 1354 57369
rect 1410 57313 1478 57369
rect 1534 57313 1602 57369
rect 1658 57313 1726 57369
rect 1782 57313 1850 57369
rect 1906 57313 2000 57369
rect 0 57200 2000 57313
rect 0 56889 2000 57000
rect 0 56833 114 56889
rect 170 56833 238 56889
rect 294 56833 362 56889
rect 418 56833 486 56889
rect 542 56833 610 56889
rect 666 56833 734 56889
rect 790 56833 858 56889
rect 914 56833 982 56889
rect 1038 56833 1106 56889
rect 1162 56833 1230 56889
rect 1286 56833 1354 56889
rect 1410 56833 1478 56889
rect 1534 56833 1602 56889
rect 1658 56833 1726 56889
rect 1782 56833 1850 56889
rect 1906 56833 2000 56889
rect 0 56765 2000 56833
rect 0 56709 114 56765
rect 170 56709 238 56765
rect 294 56709 362 56765
rect 418 56709 486 56765
rect 542 56709 610 56765
rect 666 56709 734 56765
rect 790 56709 858 56765
rect 914 56709 982 56765
rect 1038 56709 1106 56765
rect 1162 56709 1230 56765
rect 1286 56709 1354 56765
rect 1410 56709 1478 56765
rect 1534 56709 1602 56765
rect 1658 56709 1726 56765
rect 1782 56709 1850 56765
rect 1906 56709 2000 56765
rect 0 56641 2000 56709
rect 0 56585 114 56641
rect 170 56585 238 56641
rect 294 56585 362 56641
rect 418 56585 486 56641
rect 542 56585 610 56641
rect 666 56585 734 56641
rect 790 56585 858 56641
rect 914 56585 982 56641
rect 1038 56585 1106 56641
rect 1162 56585 1230 56641
rect 1286 56585 1354 56641
rect 1410 56585 1478 56641
rect 1534 56585 1602 56641
rect 1658 56585 1726 56641
rect 1782 56585 1850 56641
rect 1906 56585 2000 56641
rect 0 56517 2000 56585
rect 0 56461 114 56517
rect 170 56461 238 56517
rect 294 56461 362 56517
rect 418 56461 486 56517
rect 542 56461 610 56517
rect 666 56461 734 56517
rect 790 56461 858 56517
rect 914 56461 982 56517
rect 1038 56461 1106 56517
rect 1162 56461 1230 56517
rect 1286 56461 1354 56517
rect 1410 56461 1478 56517
rect 1534 56461 1602 56517
rect 1658 56461 1726 56517
rect 1782 56461 1850 56517
rect 1906 56461 2000 56517
rect 0 56393 2000 56461
rect 0 56337 114 56393
rect 170 56337 238 56393
rect 294 56337 362 56393
rect 418 56337 486 56393
rect 542 56337 610 56393
rect 666 56337 734 56393
rect 790 56337 858 56393
rect 914 56337 982 56393
rect 1038 56337 1106 56393
rect 1162 56337 1230 56393
rect 1286 56337 1354 56393
rect 1410 56337 1478 56393
rect 1534 56337 1602 56393
rect 1658 56337 1726 56393
rect 1782 56337 1850 56393
rect 1906 56337 2000 56393
rect 0 56269 2000 56337
rect 0 56213 114 56269
rect 170 56213 238 56269
rect 294 56213 362 56269
rect 418 56213 486 56269
rect 542 56213 610 56269
rect 666 56213 734 56269
rect 790 56213 858 56269
rect 914 56213 982 56269
rect 1038 56213 1106 56269
rect 1162 56213 1230 56269
rect 1286 56213 1354 56269
rect 1410 56213 1478 56269
rect 1534 56213 1602 56269
rect 1658 56213 1726 56269
rect 1782 56213 1850 56269
rect 1906 56213 2000 56269
rect 0 56145 2000 56213
rect 0 56089 114 56145
rect 170 56089 238 56145
rect 294 56089 362 56145
rect 418 56089 486 56145
rect 542 56089 610 56145
rect 666 56089 734 56145
rect 790 56089 858 56145
rect 914 56089 982 56145
rect 1038 56089 1106 56145
rect 1162 56089 1230 56145
rect 1286 56089 1354 56145
rect 1410 56089 1478 56145
rect 1534 56089 1602 56145
rect 1658 56089 1726 56145
rect 1782 56089 1850 56145
rect 1906 56089 2000 56145
rect 0 56021 2000 56089
rect 0 55965 114 56021
rect 170 55965 238 56021
rect 294 55965 362 56021
rect 418 55965 486 56021
rect 542 55965 610 56021
rect 666 55965 734 56021
rect 790 55965 858 56021
rect 914 55965 982 56021
rect 1038 55965 1106 56021
rect 1162 55965 1230 56021
rect 1286 55965 1354 56021
rect 1410 55965 1478 56021
rect 1534 55965 1602 56021
rect 1658 55965 1726 56021
rect 1782 55965 1850 56021
rect 1906 55965 2000 56021
rect 0 55897 2000 55965
rect 0 55841 114 55897
rect 170 55841 238 55897
rect 294 55841 362 55897
rect 418 55841 486 55897
rect 542 55841 610 55897
rect 666 55841 734 55897
rect 790 55841 858 55897
rect 914 55841 982 55897
rect 1038 55841 1106 55897
rect 1162 55841 1230 55897
rect 1286 55841 1354 55897
rect 1410 55841 1478 55897
rect 1534 55841 1602 55897
rect 1658 55841 1726 55897
rect 1782 55841 1850 55897
rect 1906 55841 2000 55897
rect 0 55773 2000 55841
rect 0 55717 114 55773
rect 170 55717 238 55773
rect 294 55717 362 55773
rect 418 55717 486 55773
rect 542 55717 610 55773
rect 666 55717 734 55773
rect 790 55717 858 55773
rect 914 55717 982 55773
rect 1038 55717 1106 55773
rect 1162 55717 1230 55773
rect 1286 55717 1354 55773
rect 1410 55717 1478 55773
rect 1534 55717 1602 55773
rect 1658 55717 1726 55773
rect 1782 55717 1850 55773
rect 1906 55717 2000 55773
rect 0 55600 2000 55717
rect 0 55280 2000 55400
rect 0 55224 114 55280
rect 170 55224 238 55280
rect 294 55224 362 55280
rect 418 55224 486 55280
rect 542 55224 610 55280
rect 666 55224 734 55280
rect 790 55224 858 55280
rect 914 55224 982 55280
rect 1038 55224 1106 55280
rect 1162 55224 1230 55280
rect 1286 55224 1354 55280
rect 1410 55224 1478 55280
rect 1534 55224 1602 55280
rect 1658 55224 1726 55280
rect 1782 55224 1850 55280
rect 1906 55224 2000 55280
rect 0 55156 2000 55224
rect 0 55100 114 55156
rect 170 55100 238 55156
rect 294 55100 362 55156
rect 418 55100 486 55156
rect 542 55100 610 55156
rect 666 55100 734 55156
rect 790 55100 858 55156
rect 914 55100 982 55156
rect 1038 55100 1106 55156
rect 1162 55100 1230 55156
rect 1286 55100 1354 55156
rect 1410 55100 1478 55156
rect 1534 55100 1602 55156
rect 1658 55100 1726 55156
rect 1782 55100 1850 55156
rect 1906 55100 2000 55156
rect 0 55032 2000 55100
rect 0 54976 114 55032
rect 170 54976 238 55032
rect 294 54976 362 55032
rect 418 54976 486 55032
rect 542 54976 610 55032
rect 666 54976 734 55032
rect 790 54976 858 55032
rect 914 54976 982 55032
rect 1038 54976 1106 55032
rect 1162 54976 1230 55032
rect 1286 54976 1354 55032
rect 1410 54976 1478 55032
rect 1534 54976 1602 55032
rect 1658 54976 1726 55032
rect 1782 54976 1850 55032
rect 1906 54976 2000 55032
rect 0 54908 2000 54976
rect 0 54852 114 54908
rect 170 54852 238 54908
rect 294 54852 362 54908
rect 418 54852 486 54908
rect 542 54852 610 54908
rect 666 54852 734 54908
rect 790 54852 858 54908
rect 914 54852 982 54908
rect 1038 54852 1106 54908
rect 1162 54852 1230 54908
rect 1286 54852 1354 54908
rect 1410 54852 1478 54908
rect 1534 54852 1602 54908
rect 1658 54852 1726 54908
rect 1782 54852 1850 54908
rect 1906 54852 2000 54908
rect 0 54784 2000 54852
rect 0 54728 114 54784
rect 170 54728 238 54784
rect 294 54728 362 54784
rect 418 54728 486 54784
rect 542 54728 610 54784
rect 666 54728 734 54784
rect 790 54728 858 54784
rect 914 54728 982 54784
rect 1038 54728 1106 54784
rect 1162 54728 1230 54784
rect 1286 54728 1354 54784
rect 1410 54728 1478 54784
rect 1534 54728 1602 54784
rect 1658 54728 1726 54784
rect 1782 54728 1850 54784
rect 1906 54728 2000 54784
rect 0 54660 2000 54728
rect 0 54604 114 54660
rect 170 54604 238 54660
rect 294 54604 362 54660
rect 418 54604 486 54660
rect 542 54604 610 54660
rect 666 54604 734 54660
rect 790 54604 858 54660
rect 914 54604 982 54660
rect 1038 54604 1106 54660
rect 1162 54604 1230 54660
rect 1286 54604 1354 54660
rect 1410 54604 1478 54660
rect 1534 54604 1602 54660
rect 1658 54604 1726 54660
rect 1782 54604 1850 54660
rect 1906 54604 2000 54660
rect 0 54536 2000 54604
rect 0 54480 114 54536
rect 170 54480 238 54536
rect 294 54480 362 54536
rect 418 54480 486 54536
rect 542 54480 610 54536
rect 666 54480 734 54536
rect 790 54480 858 54536
rect 914 54480 982 54536
rect 1038 54480 1106 54536
rect 1162 54480 1230 54536
rect 1286 54480 1354 54536
rect 1410 54480 1478 54536
rect 1534 54480 1602 54536
rect 1658 54480 1726 54536
rect 1782 54480 1850 54536
rect 1906 54480 2000 54536
rect 0 54412 2000 54480
rect 0 54356 114 54412
rect 170 54356 238 54412
rect 294 54356 362 54412
rect 418 54356 486 54412
rect 542 54356 610 54412
rect 666 54356 734 54412
rect 790 54356 858 54412
rect 914 54356 982 54412
rect 1038 54356 1106 54412
rect 1162 54356 1230 54412
rect 1286 54356 1354 54412
rect 1410 54356 1478 54412
rect 1534 54356 1602 54412
rect 1658 54356 1726 54412
rect 1782 54356 1850 54412
rect 1906 54356 2000 54412
rect 0 54288 2000 54356
rect 0 54232 114 54288
rect 170 54232 238 54288
rect 294 54232 362 54288
rect 418 54232 486 54288
rect 542 54232 610 54288
rect 666 54232 734 54288
rect 790 54232 858 54288
rect 914 54232 982 54288
rect 1038 54232 1106 54288
rect 1162 54232 1230 54288
rect 1286 54232 1354 54288
rect 1410 54232 1478 54288
rect 1534 54232 1602 54288
rect 1658 54232 1726 54288
rect 1782 54232 1850 54288
rect 1906 54232 2000 54288
rect 0 54164 2000 54232
rect 0 54108 114 54164
rect 170 54108 238 54164
rect 294 54108 362 54164
rect 418 54108 486 54164
rect 542 54108 610 54164
rect 666 54108 734 54164
rect 790 54108 858 54164
rect 914 54108 982 54164
rect 1038 54108 1106 54164
rect 1162 54108 1230 54164
rect 1286 54108 1354 54164
rect 1410 54108 1478 54164
rect 1534 54108 1602 54164
rect 1658 54108 1726 54164
rect 1782 54108 1850 54164
rect 1906 54108 2000 54164
rect 0 54000 2000 54108
rect 0 53707 2000 53800
rect 0 53651 114 53707
rect 170 53651 238 53707
rect 294 53651 362 53707
rect 418 53651 486 53707
rect 542 53651 610 53707
rect 666 53651 734 53707
rect 790 53651 858 53707
rect 914 53651 982 53707
rect 1038 53651 1106 53707
rect 1162 53651 1230 53707
rect 1286 53651 1354 53707
rect 1410 53651 1478 53707
rect 1534 53651 1602 53707
rect 1658 53651 1726 53707
rect 1782 53651 1850 53707
rect 1906 53651 2000 53707
rect 0 53583 2000 53651
rect 0 53527 114 53583
rect 170 53527 238 53583
rect 294 53527 362 53583
rect 418 53527 486 53583
rect 542 53527 610 53583
rect 666 53527 734 53583
rect 790 53527 858 53583
rect 914 53527 982 53583
rect 1038 53527 1106 53583
rect 1162 53527 1230 53583
rect 1286 53527 1354 53583
rect 1410 53527 1478 53583
rect 1534 53527 1602 53583
rect 1658 53527 1726 53583
rect 1782 53527 1850 53583
rect 1906 53527 2000 53583
rect 0 53459 2000 53527
rect 0 53403 114 53459
rect 170 53403 238 53459
rect 294 53403 362 53459
rect 418 53403 486 53459
rect 542 53403 610 53459
rect 666 53403 734 53459
rect 790 53403 858 53459
rect 914 53403 982 53459
rect 1038 53403 1106 53459
rect 1162 53403 1230 53459
rect 1286 53403 1354 53459
rect 1410 53403 1478 53459
rect 1534 53403 1602 53459
rect 1658 53403 1726 53459
rect 1782 53403 1850 53459
rect 1906 53403 2000 53459
rect 0 53335 2000 53403
rect 0 53279 114 53335
rect 170 53279 238 53335
rect 294 53279 362 53335
rect 418 53279 486 53335
rect 542 53279 610 53335
rect 666 53279 734 53335
rect 790 53279 858 53335
rect 914 53279 982 53335
rect 1038 53279 1106 53335
rect 1162 53279 1230 53335
rect 1286 53279 1354 53335
rect 1410 53279 1478 53335
rect 1534 53279 1602 53335
rect 1658 53279 1726 53335
rect 1782 53279 1850 53335
rect 1906 53279 2000 53335
rect 0 53211 2000 53279
rect 0 53155 114 53211
rect 170 53155 238 53211
rect 294 53155 362 53211
rect 418 53155 486 53211
rect 542 53155 610 53211
rect 666 53155 734 53211
rect 790 53155 858 53211
rect 914 53155 982 53211
rect 1038 53155 1106 53211
rect 1162 53155 1230 53211
rect 1286 53155 1354 53211
rect 1410 53155 1478 53211
rect 1534 53155 1602 53211
rect 1658 53155 1726 53211
rect 1782 53155 1850 53211
rect 1906 53155 2000 53211
rect 0 53087 2000 53155
rect 0 53031 114 53087
rect 170 53031 238 53087
rect 294 53031 362 53087
rect 418 53031 486 53087
rect 542 53031 610 53087
rect 666 53031 734 53087
rect 790 53031 858 53087
rect 914 53031 982 53087
rect 1038 53031 1106 53087
rect 1162 53031 1230 53087
rect 1286 53031 1354 53087
rect 1410 53031 1478 53087
rect 1534 53031 1602 53087
rect 1658 53031 1726 53087
rect 1782 53031 1850 53087
rect 1906 53031 2000 53087
rect 0 52963 2000 53031
rect 0 52907 114 52963
rect 170 52907 238 52963
rect 294 52907 362 52963
rect 418 52907 486 52963
rect 542 52907 610 52963
rect 666 52907 734 52963
rect 790 52907 858 52963
rect 914 52907 982 52963
rect 1038 52907 1106 52963
rect 1162 52907 1230 52963
rect 1286 52907 1354 52963
rect 1410 52907 1478 52963
rect 1534 52907 1602 52963
rect 1658 52907 1726 52963
rect 1782 52907 1850 52963
rect 1906 52907 2000 52963
rect 0 52839 2000 52907
rect 0 52783 114 52839
rect 170 52783 238 52839
rect 294 52783 362 52839
rect 418 52783 486 52839
rect 542 52783 610 52839
rect 666 52783 734 52839
rect 790 52783 858 52839
rect 914 52783 982 52839
rect 1038 52783 1106 52839
rect 1162 52783 1230 52839
rect 1286 52783 1354 52839
rect 1410 52783 1478 52839
rect 1534 52783 1602 52839
rect 1658 52783 1726 52839
rect 1782 52783 1850 52839
rect 1906 52783 2000 52839
rect 0 52715 2000 52783
rect 0 52659 114 52715
rect 170 52659 238 52715
rect 294 52659 362 52715
rect 418 52659 486 52715
rect 542 52659 610 52715
rect 666 52659 734 52715
rect 790 52659 858 52715
rect 914 52659 982 52715
rect 1038 52659 1106 52715
rect 1162 52659 1230 52715
rect 1286 52659 1354 52715
rect 1410 52659 1478 52715
rect 1534 52659 1602 52715
rect 1658 52659 1726 52715
rect 1782 52659 1850 52715
rect 1906 52659 2000 52715
rect 0 52591 2000 52659
rect 0 52535 114 52591
rect 170 52535 238 52591
rect 294 52535 362 52591
rect 418 52535 486 52591
rect 542 52535 610 52591
rect 666 52535 734 52591
rect 790 52535 858 52591
rect 914 52535 982 52591
rect 1038 52535 1106 52591
rect 1162 52535 1230 52591
rect 1286 52535 1354 52591
rect 1410 52535 1478 52591
rect 1534 52535 1602 52591
rect 1658 52535 1726 52591
rect 1782 52535 1850 52591
rect 1906 52535 2000 52591
rect 0 52400 2000 52535
rect 0 52100 2000 52200
rect 0 52044 114 52100
rect 170 52044 238 52100
rect 294 52044 362 52100
rect 418 52044 486 52100
rect 542 52044 610 52100
rect 666 52044 734 52100
rect 790 52044 858 52100
rect 914 52044 982 52100
rect 1038 52044 1106 52100
rect 1162 52044 1230 52100
rect 1286 52044 1354 52100
rect 1410 52044 1478 52100
rect 1534 52044 1602 52100
rect 1658 52044 1726 52100
rect 1782 52044 1850 52100
rect 1906 52044 2000 52100
rect 0 51976 2000 52044
rect 0 51920 114 51976
rect 170 51920 238 51976
rect 294 51920 362 51976
rect 418 51920 486 51976
rect 542 51920 610 51976
rect 666 51920 734 51976
rect 790 51920 858 51976
rect 914 51920 982 51976
rect 1038 51920 1106 51976
rect 1162 51920 1230 51976
rect 1286 51920 1354 51976
rect 1410 51920 1478 51976
rect 1534 51920 1602 51976
rect 1658 51920 1726 51976
rect 1782 51920 1850 51976
rect 1906 51920 2000 51976
rect 0 51852 2000 51920
rect 0 51796 114 51852
rect 170 51796 238 51852
rect 294 51796 362 51852
rect 418 51796 486 51852
rect 542 51796 610 51852
rect 666 51796 734 51852
rect 790 51796 858 51852
rect 914 51796 982 51852
rect 1038 51796 1106 51852
rect 1162 51796 1230 51852
rect 1286 51796 1354 51852
rect 1410 51796 1478 51852
rect 1534 51796 1602 51852
rect 1658 51796 1726 51852
rect 1782 51796 1850 51852
rect 1906 51796 2000 51852
rect 0 51728 2000 51796
rect 0 51672 114 51728
rect 170 51672 238 51728
rect 294 51672 362 51728
rect 418 51672 486 51728
rect 542 51672 610 51728
rect 666 51672 734 51728
rect 790 51672 858 51728
rect 914 51672 982 51728
rect 1038 51672 1106 51728
rect 1162 51672 1230 51728
rect 1286 51672 1354 51728
rect 1410 51672 1478 51728
rect 1534 51672 1602 51728
rect 1658 51672 1726 51728
rect 1782 51672 1850 51728
rect 1906 51672 2000 51728
rect 0 51604 2000 51672
rect 0 51548 114 51604
rect 170 51548 238 51604
rect 294 51548 362 51604
rect 418 51548 486 51604
rect 542 51548 610 51604
rect 666 51548 734 51604
rect 790 51548 858 51604
rect 914 51548 982 51604
rect 1038 51548 1106 51604
rect 1162 51548 1230 51604
rect 1286 51548 1354 51604
rect 1410 51548 1478 51604
rect 1534 51548 1602 51604
rect 1658 51548 1726 51604
rect 1782 51548 1850 51604
rect 1906 51548 2000 51604
rect 0 51480 2000 51548
rect 0 51424 114 51480
rect 170 51424 238 51480
rect 294 51424 362 51480
rect 418 51424 486 51480
rect 542 51424 610 51480
rect 666 51424 734 51480
rect 790 51424 858 51480
rect 914 51424 982 51480
rect 1038 51424 1106 51480
rect 1162 51424 1230 51480
rect 1286 51424 1354 51480
rect 1410 51424 1478 51480
rect 1534 51424 1602 51480
rect 1658 51424 1726 51480
rect 1782 51424 1850 51480
rect 1906 51424 2000 51480
rect 0 51356 2000 51424
rect 0 51300 114 51356
rect 170 51300 238 51356
rect 294 51300 362 51356
rect 418 51300 486 51356
rect 542 51300 610 51356
rect 666 51300 734 51356
rect 790 51300 858 51356
rect 914 51300 982 51356
rect 1038 51300 1106 51356
rect 1162 51300 1230 51356
rect 1286 51300 1354 51356
rect 1410 51300 1478 51356
rect 1534 51300 1602 51356
rect 1658 51300 1726 51356
rect 1782 51300 1850 51356
rect 1906 51300 2000 51356
rect 0 51232 2000 51300
rect 0 51176 114 51232
rect 170 51176 238 51232
rect 294 51176 362 51232
rect 418 51176 486 51232
rect 542 51176 610 51232
rect 666 51176 734 51232
rect 790 51176 858 51232
rect 914 51176 982 51232
rect 1038 51176 1106 51232
rect 1162 51176 1230 51232
rect 1286 51176 1354 51232
rect 1410 51176 1478 51232
rect 1534 51176 1602 51232
rect 1658 51176 1726 51232
rect 1782 51176 1850 51232
rect 1906 51176 2000 51232
rect 0 51108 2000 51176
rect 0 51052 114 51108
rect 170 51052 238 51108
rect 294 51052 362 51108
rect 418 51052 486 51108
rect 542 51052 610 51108
rect 666 51052 734 51108
rect 790 51052 858 51108
rect 914 51052 982 51108
rect 1038 51052 1106 51108
rect 1162 51052 1230 51108
rect 1286 51052 1354 51108
rect 1410 51052 1478 51108
rect 1534 51052 1602 51108
rect 1658 51052 1726 51108
rect 1782 51052 1850 51108
rect 1906 51052 2000 51108
rect 0 50984 2000 51052
rect 0 50928 114 50984
rect 170 50928 238 50984
rect 294 50928 362 50984
rect 418 50928 486 50984
rect 542 50928 610 50984
rect 666 50928 734 50984
rect 790 50928 858 50984
rect 914 50928 982 50984
rect 1038 50928 1106 50984
rect 1162 50928 1230 50984
rect 1286 50928 1354 50984
rect 1410 50928 1478 50984
rect 1534 50928 1602 50984
rect 1658 50928 1726 50984
rect 1782 50928 1850 50984
rect 1906 50928 2000 50984
rect 0 50800 2000 50928
rect 0 50480 2000 50600
rect 0 50424 114 50480
rect 170 50424 238 50480
rect 294 50424 362 50480
rect 418 50424 486 50480
rect 542 50424 610 50480
rect 666 50424 734 50480
rect 790 50424 858 50480
rect 914 50424 982 50480
rect 1038 50424 1106 50480
rect 1162 50424 1230 50480
rect 1286 50424 1354 50480
rect 1410 50424 1478 50480
rect 1534 50424 1602 50480
rect 1658 50424 1726 50480
rect 1782 50424 1850 50480
rect 1906 50424 2000 50480
rect 0 50356 2000 50424
rect 0 50300 114 50356
rect 170 50300 238 50356
rect 294 50300 362 50356
rect 418 50300 486 50356
rect 542 50300 610 50356
rect 666 50300 734 50356
rect 790 50300 858 50356
rect 914 50300 982 50356
rect 1038 50300 1106 50356
rect 1162 50300 1230 50356
rect 1286 50300 1354 50356
rect 1410 50300 1478 50356
rect 1534 50300 1602 50356
rect 1658 50300 1726 50356
rect 1782 50300 1850 50356
rect 1906 50300 2000 50356
rect 0 50232 2000 50300
rect 0 50176 114 50232
rect 170 50176 238 50232
rect 294 50176 362 50232
rect 418 50176 486 50232
rect 542 50176 610 50232
rect 666 50176 734 50232
rect 790 50176 858 50232
rect 914 50176 982 50232
rect 1038 50176 1106 50232
rect 1162 50176 1230 50232
rect 1286 50176 1354 50232
rect 1410 50176 1478 50232
rect 1534 50176 1602 50232
rect 1658 50176 1726 50232
rect 1782 50176 1850 50232
rect 1906 50176 2000 50232
rect 0 50108 2000 50176
rect 0 50052 114 50108
rect 170 50052 238 50108
rect 294 50052 362 50108
rect 418 50052 486 50108
rect 542 50052 610 50108
rect 666 50052 734 50108
rect 790 50052 858 50108
rect 914 50052 982 50108
rect 1038 50052 1106 50108
rect 1162 50052 1230 50108
rect 1286 50052 1354 50108
rect 1410 50052 1478 50108
rect 1534 50052 1602 50108
rect 1658 50052 1726 50108
rect 1782 50052 1850 50108
rect 1906 50052 2000 50108
rect 0 49984 2000 50052
rect 0 49928 114 49984
rect 170 49928 238 49984
rect 294 49928 362 49984
rect 418 49928 486 49984
rect 542 49928 610 49984
rect 666 49928 734 49984
rect 790 49928 858 49984
rect 914 49928 982 49984
rect 1038 49928 1106 49984
rect 1162 49928 1230 49984
rect 1286 49928 1354 49984
rect 1410 49928 1478 49984
rect 1534 49928 1602 49984
rect 1658 49928 1726 49984
rect 1782 49928 1850 49984
rect 1906 49928 2000 49984
rect 0 49860 2000 49928
rect 0 49804 114 49860
rect 170 49804 238 49860
rect 294 49804 362 49860
rect 418 49804 486 49860
rect 542 49804 610 49860
rect 666 49804 734 49860
rect 790 49804 858 49860
rect 914 49804 982 49860
rect 1038 49804 1106 49860
rect 1162 49804 1230 49860
rect 1286 49804 1354 49860
rect 1410 49804 1478 49860
rect 1534 49804 1602 49860
rect 1658 49804 1726 49860
rect 1782 49804 1850 49860
rect 1906 49804 2000 49860
rect 0 49736 2000 49804
rect 0 49680 114 49736
rect 170 49680 238 49736
rect 294 49680 362 49736
rect 418 49680 486 49736
rect 542 49680 610 49736
rect 666 49680 734 49736
rect 790 49680 858 49736
rect 914 49680 982 49736
rect 1038 49680 1106 49736
rect 1162 49680 1230 49736
rect 1286 49680 1354 49736
rect 1410 49680 1478 49736
rect 1534 49680 1602 49736
rect 1658 49680 1726 49736
rect 1782 49680 1850 49736
rect 1906 49680 2000 49736
rect 0 49612 2000 49680
rect 0 49556 114 49612
rect 170 49556 238 49612
rect 294 49556 362 49612
rect 418 49556 486 49612
rect 542 49556 610 49612
rect 666 49556 734 49612
rect 790 49556 858 49612
rect 914 49556 982 49612
rect 1038 49556 1106 49612
rect 1162 49556 1230 49612
rect 1286 49556 1354 49612
rect 1410 49556 1478 49612
rect 1534 49556 1602 49612
rect 1658 49556 1726 49612
rect 1782 49556 1850 49612
rect 1906 49556 2000 49612
rect 0 49488 2000 49556
rect 0 49432 114 49488
rect 170 49432 238 49488
rect 294 49432 362 49488
rect 418 49432 486 49488
rect 542 49432 610 49488
rect 666 49432 734 49488
rect 790 49432 858 49488
rect 914 49432 982 49488
rect 1038 49432 1106 49488
rect 1162 49432 1230 49488
rect 1286 49432 1354 49488
rect 1410 49432 1478 49488
rect 1534 49432 1602 49488
rect 1658 49432 1726 49488
rect 1782 49432 1850 49488
rect 1906 49432 2000 49488
rect 0 49364 2000 49432
rect 0 49308 114 49364
rect 170 49308 238 49364
rect 294 49308 362 49364
rect 418 49308 486 49364
rect 542 49308 610 49364
rect 666 49308 734 49364
rect 790 49308 858 49364
rect 914 49308 982 49364
rect 1038 49308 1106 49364
rect 1162 49308 1230 49364
rect 1286 49308 1354 49364
rect 1410 49308 1478 49364
rect 1534 49308 1602 49364
rect 1658 49308 1726 49364
rect 1782 49308 1850 49364
rect 1906 49308 2000 49364
rect 0 49200 2000 49308
rect 0 48841 2000 49000
rect 0 48785 114 48841
rect 170 48785 238 48841
rect 294 48785 362 48841
rect 418 48785 486 48841
rect 542 48785 610 48841
rect 666 48785 734 48841
rect 790 48785 858 48841
rect 914 48785 982 48841
rect 1038 48785 1106 48841
rect 1162 48785 1230 48841
rect 1286 48785 1354 48841
rect 1410 48785 1478 48841
rect 1534 48785 1602 48841
rect 1658 48785 1726 48841
rect 1782 48785 1850 48841
rect 1906 48785 2000 48841
rect 0 48717 2000 48785
rect 0 48661 114 48717
rect 170 48661 238 48717
rect 294 48661 362 48717
rect 418 48661 486 48717
rect 542 48661 610 48717
rect 666 48661 734 48717
rect 790 48661 858 48717
rect 914 48661 982 48717
rect 1038 48661 1106 48717
rect 1162 48661 1230 48717
rect 1286 48661 1354 48717
rect 1410 48661 1478 48717
rect 1534 48661 1602 48717
rect 1658 48661 1726 48717
rect 1782 48661 1850 48717
rect 1906 48661 2000 48717
rect 0 48593 2000 48661
rect 0 48537 114 48593
rect 170 48537 238 48593
rect 294 48537 362 48593
rect 418 48537 486 48593
rect 542 48537 610 48593
rect 666 48537 734 48593
rect 790 48537 858 48593
rect 914 48537 982 48593
rect 1038 48537 1106 48593
rect 1162 48537 1230 48593
rect 1286 48537 1354 48593
rect 1410 48537 1478 48593
rect 1534 48537 1602 48593
rect 1658 48537 1726 48593
rect 1782 48537 1850 48593
rect 1906 48537 2000 48593
rect 0 48469 2000 48537
rect 0 48413 114 48469
rect 170 48413 238 48469
rect 294 48413 362 48469
rect 418 48413 486 48469
rect 542 48413 610 48469
rect 666 48413 734 48469
rect 790 48413 858 48469
rect 914 48413 982 48469
rect 1038 48413 1106 48469
rect 1162 48413 1230 48469
rect 1286 48413 1354 48469
rect 1410 48413 1478 48469
rect 1534 48413 1602 48469
rect 1658 48413 1726 48469
rect 1782 48413 1850 48469
rect 1906 48413 2000 48469
rect 0 48345 2000 48413
rect 0 48289 114 48345
rect 170 48289 238 48345
rect 294 48289 362 48345
rect 418 48289 486 48345
rect 542 48289 610 48345
rect 666 48289 734 48345
rect 790 48289 858 48345
rect 914 48289 982 48345
rect 1038 48289 1106 48345
rect 1162 48289 1230 48345
rect 1286 48289 1354 48345
rect 1410 48289 1478 48345
rect 1534 48289 1602 48345
rect 1658 48289 1726 48345
rect 1782 48289 1850 48345
rect 1906 48289 2000 48345
rect 0 48221 2000 48289
rect 0 48165 114 48221
rect 170 48165 238 48221
rect 294 48165 362 48221
rect 418 48165 486 48221
rect 542 48165 610 48221
rect 666 48165 734 48221
rect 790 48165 858 48221
rect 914 48165 982 48221
rect 1038 48165 1106 48221
rect 1162 48165 1230 48221
rect 1286 48165 1354 48221
rect 1410 48165 1478 48221
rect 1534 48165 1602 48221
rect 1658 48165 1726 48221
rect 1782 48165 1850 48221
rect 1906 48165 2000 48221
rect 0 48097 2000 48165
rect 0 48041 114 48097
rect 170 48041 238 48097
rect 294 48041 362 48097
rect 418 48041 486 48097
rect 542 48041 610 48097
rect 666 48041 734 48097
rect 790 48041 858 48097
rect 914 48041 982 48097
rect 1038 48041 1106 48097
rect 1162 48041 1230 48097
rect 1286 48041 1354 48097
rect 1410 48041 1478 48097
rect 1534 48041 1602 48097
rect 1658 48041 1726 48097
rect 1782 48041 1850 48097
rect 1906 48041 2000 48097
rect 0 47973 2000 48041
rect 0 47917 114 47973
rect 170 47917 238 47973
rect 294 47917 362 47973
rect 418 47917 486 47973
rect 542 47917 610 47973
rect 666 47917 734 47973
rect 790 47917 858 47973
rect 914 47917 982 47973
rect 1038 47917 1106 47973
rect 1162 47917 1230 47973
rect 1286 47917 1354 47973
rect 1410 47917 1478 47973
rect 1534 47917 1602 47973
rect 1658 47917 1726 47973
rect 1782 47917 1850 47973
rect 1906 47917 2000 47973
rect 0 47849 2000 47917
rect 0 47793 114 47849
rect 170 47793 238 47849
rect 294 47793 362 47849
rect 418 47793 486 47849
rect 542 47793 610 47849
rect 666 47793 734 47849
rect 790 47793 858 47849
rect 914 47793 982 47849
rect 1038 47793 1106 47849
rect 1162 47793 1230 47849
rect 1286 47793 1354 47849
rect 1410 47793 1478 47849
rect 1534 47793 1602 47849
rect 1658 47793 1726 47849
rect 1782 47793 1850 47849
rect 1906 47793 2000 47849
rect 0 47725 2000 47793
rect 0 47669 114 47725
rect 170 47669 238 47725
rect 294 47669 362 47725
rect 418 47669 486 47725
rect 542 47669 610 47725
rect 666 47669 734 47725
rect 790 47669 858 47725
rect 914 47669 982 47725
rect 1038 47669 1106 47725
rect 1162 47669 1230 47725
rect 1286 47669 1354 47725
rect 1410 47669 1478 47725
rect 1534 47669 1602 47725
rect 1658 47669 1726 47725
rect 1782 47669 1850 47725
rect 1906 47669 2000 47725
rect 0 47601 2000 47669
rect 0 47545 114 47601
rect 170 47545 238 47601
rect 294 47545 362 47601
rect 418 47545 486 47601
rect 542 47545 610 47601
rect 666 47545 734 47601
rect 790 47545 858 47601
rect 914 47545 982 47601
rect 1038 47545 1106 47601
rect 1162 47545 1230 47601
rect 1286 47545 1354 47601
rect 1410 47545 1478 47601
rect 1534 47545 1602 47601
rect 1658 47545 1726 47601
rect 1782 47545 1850 47601
rect 1906 47545 2000 47601
rect 0 47477 2000 47545
rect 0 47421 114 47477
rect 170 47421 238 47477
rect 294 47421 362 47477
rect 418 47421 486 47477
rect 542 47421 610 47477
rect 666 47421 734 47477
rect 790 47421 858 47477
rect 914 47421 982 47477
rect 1038 47421 1106 47477
rect 1162 47421 1230 47477
rect 1286 47421 1354 47477
rect 1410 47421 1478 47477
rect 1534 47421 1602 47477
rect 1658 47421 1726 47477
rect 1782 47421 1850 47477
rect 1906 47421 2000 47477
rect 0 47353 2000 47421
rect 0 47297 114 47353
rect 170 47297 238 47353
rect 294 47297 362 47353
rect 418 47297 486 47353
rect 542 47297 610 47353
rect 666 47297 734 47353
rect 790 47297 858 47353
rect 914 47297 982 47353
rect 1038 47297 1106 47353
rect 1162 47297 1230 47353
rect 1286 47297 1354 47353
rect 1410 47297 1478 47353
rect 1534 47297 1602 47353
rect 1658 47297 1726 47353
rect 1782 47297 1850 47353
rect 1906 47297 2000 47353
rect 0 47229 2000 47297
rect 0 47173 114 47229
rect 170 47173 238 47229
rect 294 47173 362 47229
rect 418 47173 486 47229
rect 542 47173 610 47229
rect 666 47173 734 47229
rect 790 47173 858 47229
rect 914 47173 982 47229
rect 1038 47173 1106 47229
rect 1162 47173 1230 47229
rect 1286 47173 1354 47229
rect 1410 47173 1478 47229
rect 1534 47173 1602 47229
rect 1658 47173 1726 47229
rect 1782 47173 1850 47229
rect 1906 47173 2000 47229
rect 0 47105 2000 47173
rect 0 47049 114 47105
rect 170 47049 238 47105
rect 294 47049 362 47105
rect 418 47049 486 47105
rect 542 47049 610 47105
rect 666 47049 734 47105
rect 790 47049 858 47105
rect 914 47049 982 47105
rect 1038 47049 1106 47105
rect 1162 47049 1230 47105
rect 1286 47049 1354 47105
rect 1410 47049 1478 47105
rect 1534 47049 1602 47105
rect 1658 47049 1726 47105
rect 1782 47049 1850 47105
rect 1906 47049 2000 47105
rect 0 46981 2000 47049
rect 0 46925 114 46981
rect 170 46925 238 46981
rect 294 46925 362 46981
rect 418 46925 486 46981
rect 542 46925 610 46981
rect 666 46925 734 46981
rect 790 46925 858 46981
rect 914 46925 982 46981
rect 1038 46925 1106 46981
rect 1162 46925 1230 46981
rect 1286 46925 1354 46981
rect 1410 46925 1478 46981
rect 1534 46925 1602 46981
rect 1658 46925 1726 46981
rect 1782 46925 1850 46981
rect 1906 46925 2000 46981
rect 0 46857 2000 46925
rect 0 46801 114 46857
rect 170 46801 238 46857
rect 294 46801 362 46857
rect 418 46801 486 46857
rect 542 46801 610 46857
rect 666 46801 734 46857
rect 790 46801 858 46857
rect 914 46801 982 46857
rect 1038 46801 1106 46857
rect 1162 46801 1230 46857
rect 1286 46801 1354 46857
rect 1410 46801 1478 46857
rect 1534 46801 1602 46857
rect 1658 46801 1726 46857
rect 1782 46801 1850 46857
rect 1906 46801 2000 46857
rect 0 46733 2000 46801
rect 0 46677 114 46733
rect 170 46677 238 46733
rect 294 46677 362 46733
rect 418 46677 486 46733
rect 542 46677 610 46733
rect 666 46677 734 46733
rect 790 46677 858 46733
rect 914 46677 982 46733
rect 1038 46677 1106 46733
rect 1162 46677 1230 46733
rect 1286 46677 1354 46733
rect 1410 46677 1478 46733
rect 1534 46677 1602 46733
rect 1658 46677 1726 46733
rect 1782 46677 1850 46733
rect 1906 46677 2000 46733
rect 0 46609 2000 46677
rect 0 46553 114 46609
rect 170 46553 238 46609
rect 294 46553 362 46609
rect 418 46553 486 46609
rect 542 46553 610 46609
rect 666 46553 734 46609
rect 790 46553 858 46609
rect 914 46553 982 46609
rect 1038 46553 1106 46609
rect 1162 46553 1230 46609
rect 1286 46553 1354 46609
rect 1410 46553 1478 46609
rect 1534 46553 1602 46609
rect 1658 46553 1726 46609
rect 1782 46553 1850 46609
rect 1906 46553 2000 46609
rect 0 46485 2000 46553
rect 0 46429 114 46485
rect 170 46429 238 46485
rect 294 46429 362 46485
rect 418 46429 486 46485
rect 542 46429 610 46485
rect 666 46429 734 46485
rect 790 46429 858 46485
rect 914 46429 982 46485
rect 1038 46429 1106 46485
rect 1162 46429 1230 46485
rect 1286 46429 1354 46485
rect 1410 46429 1478 46485
rect 1534 46429 1602 46485
rect 1658 46429 1726 46485
rect 1782 46429 1850 46485
rect 1906 46429 2000 46485
rect 0 46361 2000 46429
rect 0 46305 114 46361
rect 170 46305 238 46361
rect 294 46305 362 46361
rect 418 46305 486 46361
rect 542 46305 610 46361
rect 666 46305 734 46361
rect 790 46305 858 46361
rect 914 46305 982 46361
rect 1038 46305 1106 46361
rect 1162 46305 1230 46361
rect 1286 46305 1354 46361
rect 1410 46305 1478 46361
rect 1534 46305 1602 46361
rect 1658 46305 1726 46361
rect 1782 46305 1850 46361
rect 1906 46305 2000 46361
rect 0 46237 2000 46305
rect 0 46181 114 46237
rect 170 46181 238 46237
rect 294 46181 362 46237
rect 418 46181 486 46237
rect 542 46181 610 46237
rect 666 46181 734 46237
rect 790 46181 858 46237
rect 914 46181 982 46237
rect 1038 46181 1106 46237
rect 1162 46181 1230 46237
rect 1286 46181 1354 46237
rect 1410 46181 1478 46237
rect 1534 46181 1602 46237
rect 1658 46181 1726 46237
rect 1782 46181 1850 46237
rect 1906 46181 2000 46237
rect 0 46000 2000 46181
rect 0 45652 2000 45800
rect 0 45596 114 45652
rect 170 45596 238 45652
rect 294 45596 362 45652
rect 418 45596 486 45652
rect 542 45596 610 45652
rect 666 45596 734 45652
rect 790 45596 858 45652
rect 914 45596 982 45652
rect 1038 45596 1106 45652
rect 1162 45596 1230 45652
rect 1286 45596 1354 45652
rect 1410 45596 1478 45652
rect 1534 45596 1602 45652
rect 1658 45596 1726 45652
rect 1782 45596 1850 45652
rect 1906 45596 2000 45652
rect 0 45528 2000 45596
rect 0 45472 114 45528
rect 170 45472 238 45528
rect 294 45472 362 45528
rect 418 45472 486 45528
rect 542 45472 610 45528
rect 666 45472 734 45528
rect 790 45472 858 45528
rect 914 45472 982 45528
rect 1038 45472 1106 45528
rect 1162 45472 1230 45528
rect 1286 45472 1354 45528
rect 1410 45472 1478 45528
rect 1534 45472 1602 45528
rect 1658 45472 1726 45528
rect 1782 45472 1850 45528
rect 1906 45472 2000 45528
rect 0 45404 2000 45472
rect 0 45348 114 45404
rect 170 45348 238 45404
rect 294 45348 362 45404
rect 418 45348 486 45404
rect 542 45348 610 45404
rect 666 45348 734 45404
rect 790 45348 858 45404
rect 914 45348 982 45404
rect 1038 45348 1106 45404
rect 1162 45348 1230 45404
rect 1286 45348 1354 45404
rect 1410 45348 1478 45404
rect 1534 45348 1602 45404
rect 1658 45348 1726 45404
rect 1782 45348 1850 45404
rect 1906 45348 2000 45404
rect 0 45280 2000 45348
rect 0 45224 114 45280
rect 170 45224 238 45280
rect 294 45224 362 45280
rect 418 45224 486 45280
rect 542 45224 610 45280
rect 666 45224 734 45280
rect 790 45224 858 45280
rect 914 45224 982 45280
rect 1038 45224 1106 45280
rect 1162 45224 1230 45280
rect 1286 45224 1354 45280
rect 1410 45224 1478 45280
rect 1534 45224 1602 45280
rect 1658 45224 1726 45280
rect 1782 45224 1850 45280
rect 1906 45224 2000 45280
rect 0 45156 2000 45224
rect 0 45100 114 45156
rect 170 45100 238 45156
rect 294 45100 362 45156
rect 418 45100 486 45156
rect 542 45100 610 45156
rect 666 45100 734 45156
rect 790 45100 858 45156
rect 914 45100 982 45156
rect 1038 45100 1106 45156
rect 1162 45100 1230 45156
rect 1286 45100 1354 45156
rect 1410 45100 1478 45156
rect 1534 45100 1602 45156
rect 1658 45100 1726 45156
rect 1782 45100 1850 45156
rect 1906 45100 2000 45156
rect 0 45032 2000 45100
rect 0 44976 114 45032
rect 170 44976 238 45032
rect 294 44976 362 45032
rect 418 44976 486 45032
rect 542 44976 610 45032
rect 666 44976 734 45032
rect 790 44976 858 45032
rect 914 44976 982 45032
rect 1038 44976 1106 45032
rect 1162 44976 1230 45032
rect 1286 44976 1354 45032
rect 1410 44976 1478 45032
rect 1534 44976 1602 45032
rect 1658 44976 1726 45032
rect 1782 44976 1850 45032
rect 1906 44976 2000 45032
rect 0 44908 2000 44976
rect 0 44852 114 44908
rect 170 44852 238 44908
rect 294 44852 362 44908
rect 418 44852 486 44908
rect 542 44852 610 44908
rect 666 44852 734 44908
rect 790 44852 858 44908
rect 914 44852 982 44908
rect 1038 44852 1106 44908
rect 1162 44852 1230 44908
rect 1286 44852 1354 44908
rect 1410 44852 1478 44908
rect 1534 44852 1602 44908
rect 1658 44852 1726 44908
rect 1782 44852 1850 44908
rect 1906 44852 2000 44908
rect 0 44784 2000 44852
rect 0 44728 114 44784
rect 170 44728 238 44784
rect 294 44728 362 44784
rect 418 44728 486 44784
rect 542 44728 610 44784
rect 666 44728 734 44784
rect 790 44728 858 44784
rect 914 44728 982 44784
rect 1038 44728 1106 44784
rect 1162 44728 1230 44784
rect 1286 44728 1354 44784
rect 1410 44728 1478 44784
rect 1534 44728 1602 44784
rect 1658 44728 1726 44784
rect 1782 44728 1850 44784
rect 1906 44728 2000 44784
rect 0 44660 2000 44728
rect 0 44604 114 44660
rect 170 44604 238 44660
rect 294 44604 362 44660
rect 418 44604 486 44660
rect 542 44604 610 44660
rect 666 44604 734 44660
rect 790 44604 858 44660
rect 914 44604 982 44660
rect 1038 44604 1106 44660
rect 1162 44604 1230 44660
rect 1286 44604 1354 44660
rect 1410 44604 1478 44660
rect 1534 44604 1602 44660
rect 1658 44604 1726 44660
rect 1782 44604 1850 44660
rect 1906 44604 2000 44660
rect 0 44536 2000 44604
rect 0 44480 114 44536
rect 170 44480 238 44536
rect 294 44480 362 44536
rect 418 44480 486 44536
rect 542 44480 610 44536
rect 666 44480 734 44536
rect 790 44480 858 44536
rect 914 44480 982 44536
rect 1038 44480 1106 44536
rect 1162 44480 1230 44536
rect 1286 44480 1354 44536
rect 1410 44480 1478 44536
rect 1534 44480 1602 44536
rect 1658 44480 1726 44536
rect 1782 44480 1850 44536
rect 1906 44480 2000 44536
rect 0 44412 2000 44480
rect 0 44356 114 44412
rect 170 44356 238 44412
rect 294 44356 362 44412
rect 418 44356 486 44412
rect 542 44356 610 44412
rect 666 44356 734 44412
rect 790 44356 858 44412
rect 914 44356 982 44412
rect 1038 44356 1106 44412
rect 1162 44356 1230 44412
rect 1286 44356 1354 44412
rect 1410 44356 1478 44412
rect 1534 44356 1602 44412
rect 1658 44356 1726 44412
rect 1782 44356 1850 44412
rect 1906 44356 2000 44412
rect 0 44288 2000 44356
rect 0 44232 114 44288
rect 170 44232 238 44288
rect 294 44232 362 44288
rect 418 44232 486 44288
rect 542 44232 610 44288
rect 666 44232 734 44288
rect 790 44232 858 44288
rect 914 44232 982 44288
rect 1038 44232 1106 44288
rect 1162 44232 1230 44288
rect 1286 44232 1354 44288
rect 1410 44232 1478 44288
rect 1534 44232 1602 44288
rect 1658 44232 1726 44288
rect 1782 44232 1850 44288
rect 1906 44232 2000 44288
rect 0 44164 2000 44232
rect 0 44108 114 44164
rect 170 44108 238 44164
rect 294 44108 362 44164
rect 418 44108 486 44164
rect 542 44108 610 44164
rect 666 44108 734 44164
rect 790 44108 858 44164
rect 914 44108 982 44164
rect 1038 44108 1106 44164
rect 1162 44108 1230 44164
rect 1286 44108 1354 44164
rect 1410 44108 1478 44164
rect 1534 44108 1602 44164
rect 1658 44108 1726 44164
rect 1782 44108 1850 44164
rect 1906 44108 2000 44164
rect 0 44040 2000 44108
rect 0 43984 114 44040
rect 170 43984 238 44040
rect 294 43984 362 44040
rect 418 43984 486 44040
rect 542 43984 610 44040
rect 666 43984 734 44040
rect 790 43984 858 44040
rect 914 43984 982 44040
rect 1038 43984 1106 44040
rect 1162 43984 1230 44040
rect 1286 43984 1354 44040
rect 1410 43984 1478 44040
rect 1534 43984 1602 44040
rect 1658 43984 1726 44040
rect 1782 43984 1850 44040
rect 1906 43984 2000 44040
rect 0 43916 2000 43984
rect 0 43860 114 43916
rect 170 43860 238 43916
rect 294 43860 362 43916
rect 418 43860 486 43916
rect 542 43860 610 43916
rect 666 43860 734 43916
rect 790 43860 858 43916
rect 914 43860 982 43916
rect 1038 43860 1106 43916
rect 1162 43860 1230 43916
rect 1286 43860 1354 43916
rect 1410 43860 1478 43916
rect 1534 43860 1602 43916
rect 1658 43860 1726 43916
rect 1782 43860 1850 43916
rect 1906 43860 2000 43916
rect 0 43792 2000 43860
rect 0 43736 114 43792
rect 170 43736 238 43792
rect 294 43736 362 43792
rect 418 43736 486 43792
rect 542 43736 610 43792
rect 666 43736 734 43792
rect 790 43736 858 43792
rect 914 43736 982 43792
rect 1038 43736 1106 43792
rect 1162 43736 1230 43792
rect 1286 43736 1354 43792
rect 1410 43736 1478 43792
rect 1534 43736 1602 43792
rect 1658 43736 1726 43792
rect 1782 43736 1850 43792
rect 1906 43736 2000 43792
rect 0 43668 2000 43736
rect 0 43612 114 43668
rect 170 43612 238 43668
rect 294 43612 362 43668
rect 418 43612 486 43668
rect 542 43612 610 43668
rect 666 43612 734 43668
rect 790 43612 858 43668
rect 914 43612 982 43668
rect 1038 43612 1106 43668
rect 1162 43612 1230 43668
rect 1286 43612 1354 43668
rect 1410 43612 1478 43668
rect 1534 43612 1602 43668
rect 1658 43612 1726 43668
rect 1782 43612 1850 43668
rect 1906 43612 2000 43668
rect 0 43544 2000 43612
rect 0 43488 114 43544
rect 170 43488 238 43544
rect 294 43488 362 43544
rect 418 43488 486 43544
rect 542 43488 610 43544
rect 666 43488 734 43544
rect 790 43488 858 43544
rect 914 43488 982 43544
rect 1038 43488 1106 43544
rect 1162 43488 1230 43544
rect 1286 43488 1354 43544
rect 1410 43488 1478 43544
rect 1534 43488 1602 43544
rect 1658 43488 1726 43544
rect 1782 43488 1850 43544
rect 1906 43488 2000 43544
rect 0 43420 2000 43488
rect 0 43364 114 43420
rect 170 43364 238 43420
rect 294 43364 362 43420
rect 418 43364 486 43420
rect 542 43364 610 43420
rect 666 43364 734 43420
rect 790 43364 858 43420
rect 914 43364 982 43420
rect 1038 43364 1106 43420
rect 1162 43364 1230 43420
rect 1286 43364 1354 43420
rect 1410 43364 1478 43420
rect 1534 43364 1602 43420
rect 1658 43364 1726 43420
rect 1782 43364 1850 43420
rect 1906 43364 2000 43420
rect 0 43296 2000 43364
rect 0 43240 114 43296
rect 170 43240 238 43296
rect 294 43240 362 43296
rect 418 43240 486 43296
rect 542 43240 610 43296
rect 666 43240 734 43296
rect 790 43240 858 43296
rect 914 43240 982 43296
rect 1038 43240 1106 43296
rect 1162 43240 1230 43296
rect 1286 43240 1354 43296
rect 1410 43240 1478 43296
rect 1534 43240 1602 43296
rect 1658 43240 1726 43296
rect 1782 43240 1850 43296
rect 1906 43240 2000 43296
rect 0 43172 2000 43240
rect 0 43116 114 43172
rect 170 43116 238 43172
rect 294 43116 362 43172
rect 418 43116 486 43172
rect 542 43116 610 43172
rect 666 43116 734 43172
rect 790 43116 858 43172
rect 914 43116 982 43172
rect 1038 43116 1106 43172
rect 1162 43116 1230 43172
rect 1286 43116 1354 43172
rect 1410 43116 1478 43172
rect 1534 43116 1602 43172
rect 1658 43116 1726 43172
rect 1782 43116 1850 43172
rect 1906 43116 2000 43172
rect 0 43048 2000 43116
rect 0 42992 114 43048
rect 170 42992 238 43048
rect 294 42992 362 43048
rect 418 42992 486 43048
rect 542 42992 610 43048
rect 666 42992 734 43048
rect 790 42992 858 43048
rect 914 42992 982 43048
rect 1038 42992 1106 43048
rect 1162 42992 1230 43048
rect 1286 42992 1354 43048
rect 1410 42992 1478 43048
rect 1534 42992 1602 43048
rect 1658 42992 1726 43048
rect 1782 42992 1850 43048
rect 1906 42992 2000 43048
rect 0 42800 2000 42992
rect 0 42487 2000 42600
rect 0 42431 114 42487
rect 170 42431 238 42487
rect 294 42431 362 42487
rect 418 42431 486 42487
rect 542 42431 610 42487
rect 666 42431 734 42487
rect 790 42431 858 42487
rect 914 42431 982 42487
rect 1038 42431 1106 42487
rect 1162 42431 1230 42487
rect 1286 42431 1354 42487
rect 1410 42431 1478 42487
rect 1534 42431 1602 42487
rect 1658 42431 1726 42487
rect 1782 42431 1850 42487
rect 1906 42431 2000 42487
rect 0 42363 2000 42431
rect 0 42307 114 42363
rect 170 42307 238 42363
rect 294 42307 362 42363
rect 418 42307 486 42363
rect 542 42307 610 42363
rect 666 42307 734 42363
rect 790 42307 858 42363
rect 914 42307 982 42363
rect 1038 42307 1106 42363
rect 1162 42307 1230 42363
rect 1286 42307 1354 42363
rect 1410 42307 1478 42363
rect 1534 42307 1602 42363
rect 1658 42307 1726 42363
rect 1782 42307 1850 42363
rect 1906 42307 2000 42363
rect 0 42239 2000 42307
rect 0 42183 114 42239
rect 170 42183 238 42239
rect 294 42183 362 42239
rect 418 42183 486 42239
rect 542 42183 610 42239
rect 666 42183 734 42239
rect 790 42183 858 42239
rect 914 42183 982 42239
rect 1038 42183 1106 42239
rect 1162 42183 1230 42239
rect 1286 42183 1354 42239
rect 1410 42183 1478 42239
rect 1534 42183 1602 42239
rect 1658 42183 1726 42239
rect 1782 42183 1850 42239
rect 1906 42183 2000 42239
rect 0 42115 2000 42183
rect 0 42059 114 42115
rect 170 42059 238 42115
rect 294 42059 362 42115
rect 418 42059 486 42115
rect 542 42059 610 42115
rect 666 42059 734 42115
rect 790 42059 858 42115
rect 914 42059 982 42115
rect 1038 42059 1106 42115
rect 1162 42059 1230 42115
rect 1286 42059 1354 42115
rect 1410 42059 1478 42115
rect 1534 42059 1602 42115
rect 1658 42059 1726 42115
rect 1782 42059 1850 42115
rect 1906 42059 2000 42115
rect 0 41991 2000 42059
rect 0 41935 114 41991
rect 170 41935 238 41991
rect 294 41935 362 41991
rect 418 41935 486 41991
rect 542 41935 610 41991
rect 666 41935 734 41991
rect 790 41935 858 41991
rect 914 41935 982 41991
rect 1038 41935 1106 41991
rect 1162 41935 1230 41991
rect 1286 41935 1354 41991
rect 1410 41935 1478 41991
rect 1534 41935 1602 41991
rect 1658 41935 1726 41991
rect 1782 41935 1850 41991
rect 1906 41935 2000 41991
rect 0 41867 2000 41935
rect 0 41811 114 41867
rect 170 41811 238 41867
rect 294 41811 362 41867
rect 418 41811 486 41867
rect 542 41811 610 41867
rect 666 41811 734 41867
rect 790 41811 858 41867
rect 914 41811 982 41867
rect 1038 41811 1106 41867
rect 1162 41811 1230 41867
rect 1286 41811 1354 41867
rect 1410 41811 1478 41867
rect 1534 41811 1602 41867
rect 1658 41811 1726 41867
rect 1782 41811 1850 41867
rect 1906 41811 2000 41867
rect 0 41743 2000 41811
rect 0 41687 114 41743
rect 170 41687 238 41743
rect 294 41687 362 41743
rect 418 41687 486 41743
rect 542 41687 610 41743
rect 666 41687 734 41743
rect 790 41687 858 41743
rect 914 41687 982 41743
rect 1038 41687 1106 41743
rect 1162 41687 1230 41743
rect 1286 41687 1354 41743
rect 1410 41687 1478 41743
rect 1534 41687 1602 41743
rect 1658 41687 1726 41743
rect 1782 41687 1850 41743
rect 1906 41687 2000 41743
rect 0 41619 2000 41687
rect 0 41563 114 41619
rect 170 41563 238 41619
rect 294 41563 362 41619
rect 418 41563 486 41619
rect 542 41563 610 41619
rect 666 41563 734 41619
rect 790 41563 858 41619
rect 914 41563 982 41619
rect 1038 41563 1106 41619
rect 1162 41563 1230 41619
rect 1286 41563 1354 41619
rect 1410 41563 1478 41619
rect 1534 41563 1602 41619
rect 1658 41563 1726 41619
rect 1782 41563 1850 41619
rect 1906 41563 2000 41619
rect 0 41495 2000 41563
rect 0 41439 114 41495
rect 170 41439 238 41495
rect 294 41439 362 41495
rect 418 41439 486 41495
rect 542 41439 610 41495
rect 666 41439 734 41495
rect 790 41439 858 41495
rect 914 41439 982 41495
rect 1038 41439 1106 41495
rect 1162 41439 1230 41495
rect 1286 41439 1354 41495
rect 1410 41439 1478 41495
rect 1534 41439 1602 41495
rect 1658 41439 1726 41495
rect 1782 41439 1850 41495
rect 1906 41439 2000 41495
rect 0 41371 2000 41439
rect 0 41315 114 41371
rect 170 41315 238 41371
rect 294 41315 362 41371
rect 418 41315 486 41371
rect 542 41315 610 41371
rect 666 41315 734 41371
rect 790 41315 858 41371
rect 914 41315 982 41371
rect 1038 41315 1106 41371
rect 1162 41315 1230 41371
rect 1286 41315 1354 41371
rect 1410 41315 1478 41371
rect 1534 41315 1602 41371
rect 1658 41315 1726 41371
rect 1782 41315 1850 41371
rect 1906 41315 2000 41371
rect 0 41200 2000 41315
rect 0 40891 2000 41000
rect 0 40835 114 40891
rect 170 40835 238 40891
rect 294 40835 362 40891
rect 418 40835 486 40891
rect 542 40835 610 40891
rect 666 40835 734 40891
rect 790 40835 858 40891
rect 914 40835 982 40891
rect 1038 40835 1106 40891
rect 1162 40835 1230 40891
rect 1286 40835 1354 40891
rect 1410 40835 1478 40891
rect 1534 40835 1602 40891
rect 1658 40835 1726 40891
rect 1782 40835 1850 40891
rect 1906 40835 2000 40891
rect 0 40767 2000 40835
rect 0 40711 114 40767
rect 170 40711 238 40767
rect 294 40711 362 40767
rect 418 40711 486 40767
rect 542 40711 610 40767
rect 666 40711 734 40767
rect 790 40711 858 40767
rect 914 40711 982 40767
rect 1038 40711 1106 40767
rect 1162 40711 1230 40767
rect 1286 40711 1354 40767
rect 1410 40711 1478 40767
rect 1534 40711 1602 40767
rect 1658 40711 1726 40767
rect 1782 40711 1850 40767
rect 1906 40711 2000 40767
rect 0 40643 2000 40711
rect 0 40587 114 40643
rect 170 40587 238 40643
rect 294 40587 362 40643
rect 418 40587 486 40643
rect 542 40587 610 40643
rect 666 40587 734 40643
rect 790 40587 858 40643
rect 914 40587 982 40643
rect 1038 40587 1106 40643
rect 1162 40587 1230 40643
rect 1286 40587 1354 40643
rect 1410 40587 1478 40643
rect 1534 40587 1602 40643
rect 1658 40587 1726 40643
rect 1782 40587 1850 40643
rect 1906 40587 2000 40643
rect 0 40519 2000 40587
rect 0 40463 114 40519
rect 170 40463 238 40519
rect 294 40463 362 40519
rect 418 40463 486 40519
rect 542 40463 610 40519
rect 666 40463 734 40519
rect 790 40463 858 40519
rect 914 40463 982 40519
rect 1038 40463 1106 40519
rect 1162 40463 1230 40519
rect 1286 40463 1354 40519
rect 1410 40463 1478 40519
rect 1534 40463 1602 40519
rect 1658 40463 1726 40519
rect 1782 40463 1850 40519
rect 1906 40463 2000 40519
rect 0 40395 2000 40463
rect 0 40339 114 40395
rect 170 40339 238 40395
rect 294 40339 362 40395
rect 418 40339 486 40395
rect 542 40339 610 40395
rect 666 40339 734 40395
rect 790 40339 858 40395
rect 914 40339 982 40395
rect 1038 40339 1106 40395
rect 1162 40339 1230 40395
rect 1286 40339 1354 40395
rect 1410 40339 1478 40395
rect 1534 40339 1602 40395
rect 1658 40339 1726 40395
rect 1782 40339 1850 40395
rect 1906 40339 2000 40395
rect 0 40271 2000 40339
rect 0 40215 114 40271
rect 170 40215 238 40271
rect 294 40215 362 40271
rect 418 40215 486 40271
rect 542 40215 610 40271
rect 666 40215 734 40271
rect 790 40215 858 40271
rect 914 40215 982 40271
rect 1038 40215 1106 40271
rect 1162 40215 1230 40271
rect 1286 40215 1354 40271
rect 1410 40215 1478 40271
rect 1534 40215 1602 40271
rect 1658 40215 1726 40271
rect 1782 40215 1850 40271
rect 1906 40215 2000 40271
rect 0 40147 2000 40215
rect 0 40091 114 40147
rect 170 40091 238 40147
rect 294 40091 362 40147
rect 418 40091 486 40147
rect 542 40091 610 40147
rect 666 40091 734 40147
rect 790 40091 858 40147
rect 914 40091 982 40147
rect 1038 40091 1106 40147
rect 1162 40091 1230 40147
rect 1286 40091 1354 40147
rect 1410 40091 1478 40147
rect 1534 40091 1602 40147
rect 1658 40091 1726 40147
rect 1782 40091 1850 40147
rect 1906 40091 2000 40147
rect 0 40023 2000 40091
rect 0 39967 114 40023
rect 170 39967 238 40023
rect 294 39967 362 40023
rect 418 39967 486 40023
rect 542 39967 610 40023
rect 666 39967 734 40023
rect 790 39967 858 40023
rect 914 39967 982 40023
rect 1038 39967 1106 40023
rect 1162 39967 1230 40023
rect 1286 39967 1354 40023
rect 1410 39967 1478 40023
rect 1534 39967 1602 40023
rect 1658 39967 1726 40023
rect 1782 39967 1850 40023
rect 1906 39967 2000 40023
rect 0 39899 2000 39967
rect 0 39843 114 39899
rect 170 39843 238 39899
rect 294 39843 362 39899
rect 418 39843 486 39899
rect 542 39843 610 39899
rect 666 39843 734 39899
rect 790 39843 858 39899
rect 914 39843 982 39899
rect 1038 39843 1106 39899
rect 1162 39843 1230 39899
rect 1286 39843 1354 39899
rect 1410 39843 1478 39899
rect 1534 39843 1602 39899
rect 1658 39843 1726 39899
rect 1782 39843 1850 39899
rect 1906 39843 2000 39899
rect 0 39775 2000 39843
rect 0 39719 114 39775
rect 170 39719 238 39775
rect 294 39719 362 39775
rect 418 39719 486 39775
rect 542 39719 610 39775
rect 666 39719 734 39775
rect 790 39719 858 39775
rect 914 39719 982 39775
rect 1038 39719 1106 39775
rect 1162 39719 1230 39775
rect 1286 39719 1354 39775
rect 1410 39719 1478 39775
rect 1534 39719 1602 39775
rect 1658 39719 1726 39775
rect 1782 39719 1850 39775
rect 1906 39719 2000 39775
rect 0 39600 2000 39719
rect 0 39244 2000 39400
rect 0 39188 114 39244
rect 170 39188 238 39244
rect 294 39188 362 39244
rect 418 39188 486 39244
rect 542 39188 610 39244
rect 666 39188 734 39244
rect 790 39188 858 39244
rect 914 39188 982 39244
rect 1038 39188 1106 39244
rect 1162 39188 1230 39244
rect 1286 39188 1354 39244
rect 1410 39188 1478 39244
rect 1534 39188 1602 39244
rect 1658 39188 1726 39244
rect 1782 39188 1850 39244
rect 1906 39188 2000 39244
rect 0 39120 2000 39188
rect 0 39064 114 39120
rect 170 39064 238 39120
rect 294 39064 362 39120
rect 418 39064 486 39120
rect 542 39064 610 39120
rect 666 39064 734 39120
rect 790 39064 858 39120
rect 914 39064 982 39120
rect 1038 39064 1106 39120
rect 1162 39064 1230 39120
rect 1286 39064 1354 39120
rect 1410 39064 1478 39120
rect 1534 39064 1602 39120
rect 1658 39064 1726 39120
rect 1782 39064 1850 39120
rect 1906 39064 2000 39120
rect 0 38996 2000 39064
rect 0 38940 114 38996
rect 170 38940 238 38996
rect 294 38940 362 38996
rect 418 38940 486 38996
rect 542 38940 610 38996
rect 666 38940 734 38996
rect 790 38940 858 38996
rect 914 38940 982 38996
rect 1038 38940 1106 38996
rect 1162 38940 1230 38996
rect 1286 38940 1354 38996
rect 1410 38940 1478 38996
rect 1534 38940 1602 38996
rect 1658 38940 1726 38996
rect 1782 38940 1850 38996
rect 1906 38940 2000 38996
rect 0 38872 2000 38940
rect 0 38816 114 38872
rect 170 38816 238 38872
rect 294 38816 362 38872
rect 418 38816 486 38872
rect 542 38816 610 38872
rect 666 38816 734 38872
rect 790 38816 858 38872
rect 914 38816 982 38872
rect 1038 38816 1106 38872
rect 1162 38816 1230 38872
rect 1286 38816 1354 38872
rect 1410 38816 1478 38872
rect 1534 38816 1602 38872
rect 1658 38816 1726 38872
rect 1782 38816 1850 38872
rect 1906 38816 2000 38872
rect 0 38748 2000 38816
rect 0 38692 114 38748
rect 170 38692 238 38748
rect 294 38692 362 38748
rect 418 38692 486 38748
rect 542 38692 610 38748
rect 666 38692 734 38748
rect 790 38692 858 38748
rect 914 38692 982 38748
rect 1038 38692 1106 38748
rect 1162 38692 1230 38748
rect 1286 38692 1354 38748
rect 1410 38692 1478 38748
rect 1534 38692 1602 38748
rect 1658 38692 1726 38748
rect 1782 38692 1850 38748
rect 1906 38692 2000 38748
rect 0 38624 2000 38692
rect 0 38568 114 38624
rect 170 38568 238 38624
rect 294 38568 362 38624
rect 418 38568 486 38624
rect 542 38568 610 38624
rect 666 38568 734 38624
rect 790 38568 858 38624
rect 914 38568 982 38624
rect 1038 38568 1106 38624
rect 1162 38568 1230 38624
rect 1286 38568 1354 38624
rect 1410 38568 1478 38624
rect 1534 38568 1602 38624
rect 1658 38568 1726 38624
rect 1782 38568 1850 38624
rect 1906 38568 2000 38624
rect 0 38500 2000 38568
rect 0 38444 114 38500
rect 170 38444 238 38500
rect 294 38444 362 38500
rect 418 38444 486 38500
rect 542 38444 610 38500
rect 666 38444 734 38500
rect 790 38444 858 38500
rect 914 38444 982 38500
rect 1038 38444 1106 38500
rect 1162 38444 1230 38500
rect 1286 38444 1354 38500
rect 1410 38444 1478 38500
rect 1534 38444 1602 38500
rect 1658 38444 1726 38500
rect 1782 38444 1850 38500
rect 1906 38444 2000 38500
rect 0 38376 2000 38444
rect 0 38320 114 38376
rect 170 38320 238 38376
rect 294 38320 362 38376
rect 418 38320 486 38376
rect 542 38320 610 38376
rect 666 38320 734 38376
rect 790 38320 858 38376
rect 914 38320 982 38376
rect 1038 38320 1106 38376
rect 1162 38320 1230 38376
rect 1286 38320 1354 38376
rect 1410 38320 1478 38376
rect 1534 38320 1602 38376
rect 1658 38320 1726 38376
rect 1782 38320 1850 38376
rect 1906 38320 2000 38376
rect 0 38252 2000 38320
rect 0 38196 114 38252
rect 170 38196 238 38252
rect 294 38196 362 38252
rect 418 38196 486 38252
rect 542 38196 610 38252
rect 666 38196 734 38252
rect 790 38196 858 38252
rect 914 38196 982 38252
rect 1038 38196 1106 38252
rect 1162 38196 1230 38252
rect 1286 38196 1354 38252
rect 1410 38196 1478 38252
rect 1534 38196 1602 38252
rect 1658 38196 1726 38252
rect 1782 38196 1850 38252
rect 1906 38196 2000 38252
rect 0 38128 2000 38196
rect 0 38072 114 38128
rect 170 38072 238 38128
rect 294 38072 362 38128
rect 418 38072 486 38128
rect 542 38072 610 38128
rect 666 38072 734 38128
rect 790 38072 858 38128
rect 914 38072 982 38128
rect 1038 38072 1106 38128
rect 1162 38072 1230 38128
rect 1286 38072 1354 38128
rect 1410 38072 1478 38128
rect 1534 38072 1602 38128
rect 1658 38072 1726 38128
rect 1782 38072 1850 38128
rect 1906 38072 2000 38128
rect 0 38004 2000 38072
rect 0 37948 114 38004
rect 170 37948 238 38004
rect 294 37948 362 38004
rect 418 37948 486 38004
rect 542 37948 610 38004
rect 666 37948 734 38004
rect 790 37948 858 38004
rect 914 37948 982 38004
rect 1038 37948 1106 38004
rect 1162 37948 1230 38004
rect 1286 37948 1354 38004
rect 1410 37948 1478 38004
rect 1534 37948 1602 38004
rect 1658 37948 1726 38004
rect 1782 37948 1850 38004
rect 1906 37948 2000 38004
rect 0 37880 2000 37948
rect 0 37824 114 37880
rect 170 37824 238 37880
rect 294 37824 362 37880
rect 418 37824 486 37880
rect 542 37824 610 37880
rect 666 37824 734 37880
rect 790 37824 858 37880
rect 914 37824 982 37880
rect 1038 37824 1106 37880
rect 1162 37824 1230 37880
rect 1286 37824 1354 37880
rect 1410 37824 1478 37880
rect 1534 37824 1602 37880
rect 1658 37824 1726 37880
rect 1782 37824 1850 37880
rect 1906 37824 2000 37880
rect 0 37756 2000 37824
rect 0 37700 114 37756
rect 170 37700 238 37756
rect 294 37700 362 37756
rect 418 37700 486 37756
rect 542 37700 610 37756
rect 666 37700 734 37756
rect 790 37700 858 37756
rect 914 37700 982 37756
rect 1038 37700 1106 37756
rect 1162 37700 1230 37756
rect 1286 37700 1354 37756
rect 1410 37700 1478 37756
rect 1534 37700 1602 37756
rect 1658 37700 1726 37756
rect 1782 37700 1850 37756
rect 1906 37700 2000 37756
rect 0 37632 2000 37700
rect 0 37576 114 37632
rect 170 37576 238 37632
rect 294 37576 362 37632
rect 418 37576 486 37632
rect 542 37576 610 37632
rect 666 37576 734 37632
rect 790 37576 858 37632
rect 914 37576 982 37632
rect 1038 37576 1106 37632
rect 1162 37576 1230 37632
rect 1286 37576 1354 37632
rect 1410 37576 1478 37632
rect 1534 37576 1602 37632
rect 1658 37576 1726 37632
rect 1782 37576 1850 37632
rect 1906 37576 2000 37632
rect 0 37508 2000 37576
rect 0 37452 114 37508
rect 170 37452 238 37508
rect 294 37452 362 37508
rect 418 37452 486 37508
rect 542 37452 610 37508
rect 666 37452 734 37508
rect 790 37452 858 37508
rect 914 37452 982 37508
rect 1038 37452 1106 37508
rect 1162 37452 1230 37508
rect 1286 37452 1354 37508
rect 1410 37452 1478 37508
rect 1534 37452 1602 37508
rect 1658 37452 1726 37508
rect 1782 37452 1850 37508
rect 1906 37452 2000 37508
rect 0 37384 2000 37452
rect 0 37328 114 37384
rect 170 37328 238 37384
rect 294 37328 362 37384
rect 418 37328 486 37384
rect 542 37328 610 37384
rect 666 37328 734 37384
rect 790 37328 858 37384
rect 914 37328 982 37384
rect 1038 37328 1106 37384
rect 1162 37328 1230 37384
rect 1286 37328 1354 37384
rect 1410 37328 1478 37384
rect 1534 37328 1602 37384
rect 1658 37328 1726 37384
rect 1782 37328 1850 37384
rect 1906 37328 2000 37384
rect 0 37260 2000 37328
rect 0 37204 114 37260
rect 170 37204 238 37260
rect 294 37204 362 37260
rect 418 37204 486 37260
rect 542 37204 610 37260
rect 666 37204 734 37260
rect 790 37204 858 37260
rect 914 37204 982 37260
rect 1038 37204 1106 37260
rect 1162 37204 1230 37260
rect 1286 37204 1354 37260
rect 1410 37204 1478 37260
rect 1534 37204 1602 37260
rect 1658 37204 1726 37260
rect 1782 37204 1850 37260
rect 1906 37204 2000 37260
rect 0 37136 2000 37204
rect 0 37080 114 37136
rect 170 37080 238 37136
rect 294 37080 362 37136
rect 418 37080 486 37136
rect 542 37080 610 37136
rect 666 37080 734 37136
rect 790 37080 858 37136
rect 914 37080 982 37136
rect 1038 37080 1106 37136
rect 1162 37080 1230 37136
rect 1286 37080 1354 37136
rect 1410 37080 1478 37136
rect 1534 37080 1602 37136
rect 1658 37080 1726 37136
rect 1782 37080 1850 37136
rect 1906 37080 2000 37136
rect 0 37012 2000 37080
rect 0 36956 114 37012
rect 170 36956 238 37012
rect 294 36956 362 37012
rect 418 36956 486 37012
rect 542 36956 610 37012
rect 666 36956 734 37012
rect 790 36956 858 37012
rect 914 36956 982 37012
rect 1038 36956 1106 37012
rect 1162 36956 1230 37012
rect 1286 36956 1354 37012
rect 1410 36956 1478 37012
rect 1534 36956 1602 37012
rect 1658 36956 1726 37012
rect 1782 36956 1850 37012
rect 1906 36956 2000 37012
rect 0 36888 2000 36956
rect 0 36832 114 36888
rect 170 36832 238 36888
rect 294 36832 362 36888
rect 418 36832 486 36888
rect 542 36832 610 36888
rect 666 36832 734 36888
rect 790 36832 858 36888
rect 914 36832 982 36888
rect 1038 36832 1106 36888
rect 1162 36832 1230 36888
rect 1286 36832 1354 36888
rect 1410 36832 1478 36888
rect 1534 36832 1602 36888
rect 1658 36832 1726 36888
rect 1782 36832 1850 36888
rect 1906 36832 2000 36888
rect 0 36764 2000 36832
rect 0 36708 114 36764
rect 170 36708 238 36764
rect 294 36708 362 36764
rect 418 36708 486 36764
rect 542 36708 610 36764
rect 666 36708 734 36764
rect 790 36708 858 36764
rect 914 36708 982 36764
rect 1038 36708 1106 36764
rect 1162 36708 1230 36764
rect 1286 36708 1354 36764
rect 1410 36708 1478 36764
rect 1534 36708 1602 36764
rect 1658 36708 1726 36764
rect 1782 36708 1850 36764
rect 1906 36708 2000 36764
rect 0 36640 2000 36708
rect 0 36584 114 36640
rect 170 36584 238 36640
rect 294 36584 362 36640
rect 418 36584 486 36640
rect 542 36584 610 36640
rect 666 36584 734 36640
rect 790 36584 858 36640
rect 914 36584 982 36640
rect 1038 36584 1106 36640
rect 1162 36584 1230 36640
rect 1286 36584 1354 36640
rect 1410 36584 1478 36640
rect 1534 36584 1602 36640
rect 1658 36584 1726 36640
rect 1782 36584 1850 36640
rect 1906 36584 2000 36640
rect 0 36400 2000 36584
rect 0 36059 2000 36200
rect 0 36003 114 36059
rect 170 36003 238 36059
rect 294 36003 362 36059
rect 418 36003 486 36059
rect 542 36003 610 36059
rect 666 36003 734 36059
rect 790 36003 858 36059
rect 914 36003 982 36059
rect 1038 36003 1106 36059
rect 1162 36003 1230 36059
rect 1286 36003 1354 36059
rect 1410 36003 1478 36059
rect 1534 36003 1602 36059
rect 1658 36003 1726 36059
rect 1782 36003 1850 36059
rect 1906 36003 2000 36059
rect 0 35935 2000 36003
rect 0 35879 114 35935
rect 170 35879 238 35935
rect 294 35879 362 35935
rect 418 35879 486 35935
rect 542 35879 610 35935
rect 666 35879 734 35935
rect 790 35879 858 35935
rect 914 35879 982 35935
rect 1038 35879 1106 35935
rect 1162 35879 1230 35935
rect 1286 35879 1354 35935
rect 1410 35879 1478 35935
rect 1534 35879 1602 35935
rect 1658 35879 1726 35935
rect 1782 35879 1850 35935
rect 1906 35879 2000 35935
rect 0 35811 2000 35879
rect 0 35755 114 35811
rect 170 35755 238 35811
rect 294 35755 362 35811
rect 418 35755 486 35811
rect 542 35755 610 35811
rect 666 35755 734 35811
rect 790 35755 858 35811
rect 914 35755 982 35811
rect 1038 35755 1106 35811
rect 1162 35755 1230 35811
rect 1286 35755 1354 35811
rect 1410 35755 1478 35811
rect 1534 35755 1602 35811
rect 1658 35755 1726 35811
rect 1782 35755 1850 35811
rect 1906 35755 2000 35811
rect 0 35687 2000 35755
rect 0 35631 114 35687
rect 170 35631 238 35687
rect 294 35631 362 35687
rect 418 35631 486 35687
rect 542 35631 610 35687
rect 666 35631 734 35687
rect 790 35631 858 35687
rect 914 35631 982 35687
rect 1038 35631 1106 35687
rect 1162 35631 1230 35687
rect 1286 35631 1354 35687
rect 1410 35631 1478 35687
rect 1534 35631 1602 35687
rect 1658 35631 1726 35687
rect 1782 35631 1850 35687
rect 1906 35631 2000 35687
rect 0 35563 2000 35631
rect 0 35507 114 35563
rect 170 35507 238 35563
rect 294 35507 362 35563
rect 418 35507 486 35563
rect 542 35507 610 35563
rect 666 35507 734 35563
rect 790 35507 858 35563
rect 914 35507 982 35563
rect 1038 35507 1106 35563
rect 1162 35507 1230 35563
rect 1286 35507 1354 35563
rect 1410 35507 1478 35563
rect 1534 35507 1602 35563
rect 1658 35507 1726 35563
rect 1782 35507 1850 35563
rect 1906 35507 2000 35563
rect 0 35439 2000 35507
rect 0 35383 114 35439
rect 170 35383 238 35439
rect 294 35383 362 35439
rect 418 35383 486 35439
rect 542 35383 610 35439
rect 666 35383 734 35439
rect 790 35383 858 35439
rect 914 35383 982 35439
rect 1038 35383 1106 35439
rect 1162 35383 1230 35439
rect 1286 35383 1354 35439
rect 1410 35383 1478 35439
rect 1534 35383 1602 35439
rect 1658 35383 1726 35439
rect 1782 35383 1850 35439
rect 1906 35383 2000 35439
rect 0 35315 2000 35383
rect 0 35259 114 35315
rect 170 35259 238 35315
rect 294 35259 362 35315
rect 418 35259 486 35315
rect 542 35259 610 35315
rect 666 35259 734 35315
rect 790 35259 858 35315
rect 914 35259 982 35315
rect 1038 35259 1106 35315
rect 1162 35259 1230 35315
rect 1286 35259 1354 35315
rect 1410 35259 1478 35315
rect 1534 35259 1602 35315
rect 1658 35259 1726 35315
rect 1782 35259 1850 35315
rect 1906 35259 2000 35315
rect 0 35191 2000 35259
rect 0 35135 114 35191
rect 170 35135 238 35191
rect 294 35135 362 35191
rect 418 35135 486 35191
rect 542 35135 610 35191
rect 666 35135 734 35191
rect 790 35135 858 35191
rect 914 35135 982 35191
rect 1038 35135 1106 35191
rect 1162 35135 1230 35191
rect 1286 35135 1354 35191
rect 1410 35135 1478 35191
rect 1534 35135 1602 35191
rect 1658 35135 1726 35191
rect 1782 35135 1850 35191
rect 1906 35135 2000 35191
rect 0 35067 2000 35135
rect 0 35011 114 35067
rect 170 35011 238 35067
rect 294 35011 362 35067
rect 418 35011 486 35067
rect 542 35011 610 35067
rect 666 35011 734 35067
rect 790 35011 858 35067
rect 914 35011 982 35067
rect 1038 35011 1106 35067
rect 1162 35011 1230 35067
rect 1286 35011 1354 35067
rect 1410 35011 1478 35067
rect 1534 35011 1602 35067
rect 1658 35011 1726 35067
rect 1782 35011 1850 35067
rect 1906 35011 2000 35067
rect 0 34943 2000 35011
rect 0 34887 114 34943
rect 170 34887 238 34943
rect 294 34887 362 34943
rect 418 34887 486 34943
rect 542 34887 610 34943
rect 666 34887 734 34943
rect 790 34887 858 34943
rect 914 34887 982 34943
rect 1038 34887 1106 34943
rect 1162 34887 1230 34943
rect 1286 34887 1354 34943
rect 1410 34887 1478 34943
rect 1534 34887 1602 34943
rect 1658 34887 1726 34943
rect 1782 34887 1850 34943
rect 1906 34887 2000 34943
rect 0 34819 2000 34887
rect 0 34763 114 34819
rect 170 34763 238 34819
rect 294 34763 362 34819
rect 418 34763 486 34819
rect 542 34763 610 34819
rect 666 34763 734 34819
rect 790 34763 858 34819
rect 914 34763 982 34819
rect 1038 34763 1106 34819
rect 1162 34763 1230 34819
rect 1286 34763 1354 34819
rect 1410 34763 1478 34819
rect 1534 34763 1602 34819
rect 1658 34763 1726 34819
rect 1782 34763 1850 34819
rect 1906 34763 2000 34819
rect 0 34695 2000 34763
rect 0 34639 114 34695
rect 170 34639 238 34695
rect 294 34639 362 34695
rect 418 34639 486 34695
rect 542 34639 610 34695
rect 666 34639 734 34695
rect 790 34639 858 34695
rect 914 34639 982 34695
rect 1038 34639 1106 34695
rect 1162 34639 1230 34695
rect 1286 34639 1354 34695
rect 1410 34639 1478 34695
rect 1534 34639 1602 34695
rect 1658 34639 1726 34695
rect 1782 34639 1850 34695
rect 1906 34639 2000 34695
rect 0 34571 2000 34639
rect 0 34515 114 34571
rect 170 34515 238 34571
rect 294 34515 362 34571
rect 418 34515 486 34571
rect 542 34515 610 34571
rect 666 34515 734 34571
rect 790 34515 858 34571
rect 914 34515 982 34571
rect 1038 34515 1106 34571
rect 1162 34515 1230 34571
rect 1286 34515 1354 34571
rect 1410 34515 1478 34571
rect 1534 34515 1602 34571
rect 1658 34515 1726 34571
rect 1782 34515 1850 34571
rect 1906 34515 2000 34571
rect 0 34447 2000 34515
rect 0 34391 114 34447
rect 170 34391 238 34447
rect 294 34391 362 34447
rect 418 34391 486 34447
rect 542 34391 610 34447
rect 666 34391 734 34447
rect 790 34391 858 34447
rect 914 34391 982 34447
rect 1038 34391 1106 34447
rect 1162 34391 1230 34447
rect 1286 34391 1354 34447
rect 1410 34391 1478 34447
rect 1534 34391 1602 34447
rect 1658 34391 1726 34447
rect 1782 34391 1850 34447
rect 1906 34391 2000 34447
rect 0 34323 2000 34391
rect 0 34267 114 34323
rect 170 34267 238 34323
rect 294 34267 362 34323
rect 418 34267 486 34323
rect 542 34267 610 34323
rect 666 34267 734 34323
rect 790 34267 858 34323
rect 914 34267 982 34323
rect 1038 34267 1106 34323
rect 1162 34267 1230 34323
rect 1286 34267 1354 34323
rect 1410 34267 1478 34323
rect 1534 34267 1602 34323
rect 1658 34267 1726 34323
rect 1782 34267 1850 34323
rect 1906 34267 2000 34323
rect 0 34199 2000 34267
rect 0 34143 114 34199
rect 170 34143 238 34199
rect 294 34143 362 34199
rect 418 34143 486 34199
rect 542 34143 610 34199
rect 666 34143 734 34199
rect 790 34143 858 34199
rect 914 34143 982 34199
rect 1038 34143 1106 34199
rect 1162 34143 1230 34199
rect 1286 34143 1354 34199
rect 1410 34143 1478 34199
rect 1534 34143 1602 34199
rect 1658 34143 1726 34199
rect 1782 34143 1850 34199
rect 1906 34143 2000 34199
rect 0 34075 2000 34143
rect 0 34019 114 34075
rect 170 34019 238 34075
rect 294 34019 362 34075
rect 418 34019 486 34075
rect 542 34019 610 34075
rect 666 34019 734 34075
rect 790 34019 858 34075
rect 914 34019 982 34075
rect 1038 34019 1106 34075
rect 1162 34019 1230 34075
rect 1286 34019 1354 34075
rect 1410 34019 1478 34075
rect 1534 34019 1602 34075
rect 1658 34019 1726 34075
rect 1782 34019 1850 34075
rect 1906 34019 2000 34075
rect 0 33951 2000 34019
rect 0 33895 114 33951
rect 170 33895 238 33951
rect 294 33895 362 33951
rect 418 33895 486 33951
rect 542 33895 610 33951
rect 666 33895 734 33951
rect 790 33895 858 33951
rect 914 33895 982 33951
rect 1038 33895 1106 33951
rect 1162 33895 1230 33951
rect 1286 33895 1354 33951
rect 1410 33895 1478 33951
rect 1534 33895 1602 33951
rect 1658 33895 1726 33951
rect 1782 33895 1850 33951
rect 1906 33895 2000 33951
rect 0 33827 2000 33895
rect 0 33771 114 33827
rect 170 33771 238 33827
rect 294 33771 362 33827
rect 418 33771 486 33827
rect 542 33771 610 33827
rect 666 33771 734 33827
rect 790 33771 858 33827
rect 914 33771 982 33827
rect 1038 33771 1106 33827
rect 1162 33771 1230 33827
rect 1286 33771 1354 33827
rect 1410 33771 1478 33827
rect 1534 33771 1602 33827
rect 1658 33771 1726 33827
rect 1782 33771 1850 33827
rect 1906 33771 2000 33827
rect 0 33703 2000 33771
rect 0 33647 114 33703
rect 170 33647 238 33703
rect 294 33647 362 33703
rect 418 33647 486 33703
rect 542 33647 610 33703
rect 666 33647 734 33703
rect 790 33647 858 33703
rect 914 33647 982 33703
rect 1038 33647 1106 33703
rect 1162 33647 1230 33703
rect 1286 33647 1354 33703
rect 1410 33647 1478 33703
rect 1534 33647 1602 33703
rect 1658 33647 1726 33703
rect 1782 33647 1850 33703
rect 1906 33647 2000 33703
rect 0 33579 2000 33647
rect 0 33523 114 33579
rect 170 33523 238 33579
rect 294 33523 362 33579
rect 418 33523 486 33579
rect 542 33523 610 33579
rect 666 33523 734 33579
rect 790 33523 858 33579
rect 914 33523 982 33579
rect 1038 33523 1106 33579
rect 1162 33523 1230 33579
rect 1286 33523 1354 33579
rect 1410 33523 1478 33579
rect 1534 33523 1602 33579
rect 1658 33523 1726 33579
rect 1782 33523 1850 33579
rect 1906 33523 2000 33579
rect 0 33455 2000 33523
rect 0 33399 114 33455
rect 170 33399 238 33455
rect 294 33399 362 33455
rect 418 33399 486 33455
rect 542 33399 610 33455
rect 666 33399 734 33455
rect 790 33399 858 33455
rect 914 33399 982 33455
rect 1038 33399 1106 33455
rect 1162 33399 1230 33455
rect 1286 33399 1354 33455
rect 1410 33399 1478 33455
rect 1534 33399 1602 33455
rect 1658 33399 1726 33455
rect 1782 33399 1850 33455
rect 1906 33399 2000 33455
rect 0 33200 2000 33399
rect 0 32844 2000 33000
rect 0 32788 114 32844
rect 170 32788 238 32844
rect 294 32788 362 32844
rect 418 32788 486 32844
rect 542 32788 610 32844
rect 666 32788 734 32844
rect 790 32788 858 32844
rect 914 32788 982 32844
rect 1038 32788 1106 32844
rect 1162 32788 1230 32844
rect 1286 32788 1354 32844
rect 1410 32788 1478 32844
rect 1534 32788 1602 32844
rect 1658 32788 1726 32844
rect 1782 32788 1850 32844
rect 1906 32788 2000 32844
rect 0 32720 2000 32788
rect 0 32664 114 32720
rect 170 32664 238 32720
rect 294 32664 362 32720
rect 418 32664 486 32720
rect 542 32664 610 32720
rect 666 32664 734 32720
rect 790 32664 858 32720
rect 914 32664 982 32720
rect 1038 32664 1106 32720
rect 1162 32664 1230 32720
rect 1286 32664 1354 32720
rect 1410 32664 1478 32720
rect 1534 32664 1602 32720
rect 1658 32664 1726 32720
rect 1782 32664 1850 32720
rect 1906 32664 2000 32720
rect 0 32596 2000 32664
rect 0 32540 114 32596
rect 170 32540 238 32596
rect 294 32540 362 32596
rect 418 32540 486 32596
rect 542 32540 610 32596
rect 666 32540 734 32596
rect 790 32540 858 32596
rect 914 32540 982 32596
rect 1038 32540 1106 32596
rect 1162 32540 1230 32596
rect 1286 32540 1354 32596
rect 1410 32540 1478 32596
rect 1534 32540 1602 32596
rect 1658 32540 1726 32596
rect 1782 32540 1850 32596
rect 1906 32540 2000 32596
rect 0 32472 2000 32540
rect 0 32416 114 32472
rect 170 32416 238 32472
rect 294 32416 362 32472
rect 418 32416 486 32472
rect 542 32416 610 32472
rect 666 32416 734 32472
rect 790 32416 858 32472
rect 914 32416 982 32472
rect 1038 32416 1106 32472
rect 1162 32416 1230 32472
rect 1286 32416 1354 32472
rect 1410 32416 1478 32472
rect 1534 32416 1602 32472
rect 1658 32416 1726 32472
rect 1782 32416 1850 32472
rect 1906 32416 2000 32472
rect 0 32348 2000 32416
rect 0 32292 114 32348
rect 170 32292 238 32348
rect 294 32292 362 32348
rect 418 32292 486 32348
rect 542 32292 610 32348
rect 666 32292 734 32348
rect 790 32292 858 32348
rect 914 32292 982 32348
rect 1038 32292 1106 32348
rect 1162 32292 1230 32348
rect 1286 32292 1354 32348
rect 1410 32292 1478 32348
rect 1534 32292 1602 32348
rect 1658 32292 1726 32348
rect 1782 32292 1850 32348
rect 1906 32292 2000 32348
rect 0 32224 2000 32292
rect 0 32168 114 32224
rect 170 32168 238 32224
rect 294 32168 362 32224
rect 418 32168 486 32224
rect 542 32168 610 32224
rect 666 32168 734 32224
rect 790 32168 858 32224
rect 914 32168 982 32224
rect 1038 32168 1106 32224
rect 1162 32168 1230 32224
rect 1286 32168 1354 32224
rect 1410 32168 1478 32224
rect 1534 32168 1602 32224
rect 1658 32168 1726 32224
rect 1782 32168 1850 32224
rect 1906 32168 2000 32224
rect 0 32100 2000 32168
rect 0 32044 114 32100
rect 170 32044 238 32100
rect 294 32044 362 32100
rect 418 32044 486 32100
rect 542 32044 610 32100
rect 666 32044 734 32100
rect 790 32044 858 32100
rect 914 32044 982 32100
rect 1038 32044 1106 32100
rect 1162 32044 1230 32100
rect 1286 32044 1354 32100
rect 1410 32044 1478 32100
rect 1534 32044 1602 32100
rect 1658 32044 1726 32100
rect 1782 32044 1850 32100
rect 1906 32044 2000 32100
rect 0 31976 2000 32044
rect 0 31920 114 31976
rect 170 31920 238 31976
rect 294 31920 362 31976
rect 418 31920 486 31976
rect 542 31920 610 31976
rect 666 31920 734 31976
rect 790 31920 858 31976
rect 914 31920 982 31976
rect 1038 31920 1106 31976
rect 1162 31920 1230 31976
rect 1286 31920 1354 31976
rect 1410 31920 1478 31976
rect 1534 31920 1602 31976
rect 1658 31920 1726 31976
rect 1782 31920 1850 31976
rect 1906 31920 2000 31976
rect 0 31852 2000 31920
rect 0 31796 114 31852
rect 170 31796 238 31852
rect 294 31796 362 31852
rect 418 31796 486 31852
rect 542 31796 610 31852
rect 666 31796 734 31852
rect 790 31796 858 31852
rect 914 31796 982 31852
rect 1038 31796 1106 31852
rect 1162 31796 1230 31852
rect 1286 31796 1354 31852
rect 1410 31796 1478 31852
rect 1534 31796 1602 31852
rect 1658 31796 1726 31852
rect 1782 31796 1850 31852
rect 1906 31796 2000 31852
rect 0 31728 2000 31796
rect 0 31672 114 31728
rect 170 31672 238 31728
rect 294 31672 362 31728
rect 418 31672 486 31728
rect 542 31672 610 31728
rect 666 31672 734 31728
rect 790 31672 858 31728
rect 914 31672 982 31728
rect 1038 31672 1106 31728
rect 1162 31672 1230 31728
rect 1286 31672 1354 31728
rect 1410 31672 1478 31728
rect 1534 31672 1602 31728
rect 1658 31672 1726 31728
rect 1782 31672 1850 31728
rect 1906 31672 2000 31728
rect 0 31604 2000 31672
rect 0 31548 114 31604
rect 170 31548 238 31604
rect 294 31548 362 31604
rect 418 31548 486 31604
rect 542 31548 610 31604
rect 666 31548 734 31604
rect 790 31548 858 31604
rect 914 31548 982 31604
rect 1038 31548 1106 31604
rect 1162 31548 1230 31604
rect 1286 31548 1354 31604
rect 1410 31548 1478 31604
rect 1534 31548 1602 31604
rect 1658 31548 1726 31604
rect 1782 31548 1850 31604
rect 1906 31548 2000 31604
rect 0 31480 2000 31548
rect 0 31424 114 31480
rect 170 31424 238 31480
rect 294 31424 362 31480
rect 418 31424 486 31480
rect 542 31424 610 31480
rect 666 31424 734 31480
rect 790 31424 858 31480
rect 914 31424 982 31480
rect 1038 31424 1106 31480
rect 1162 31424 1230 31480
rect 1286 31424 1354 31480
rect 1410 31424 1478 31480
rect 1534 31424 1602 31480
rect 1658 31424 1726 31480
rect 1782 31424 1850 31480
rect 1906 31424 2000 31480
rect 0 31356 2000 31424
rect 0 31300 114 31356
rect 170 31300 238 31356
rect 294 31300 362 31356
rect 418 31300 486 31356
rect 542 31300 610 31356
rect 666 31300 734 31356
rect 790 31300 858 31356
rect 914 31300 982 31356
rect 1038 31300 1106 31356
rect 1162 31300 1230 31356
rect 1286 31300 1354 31356
rect 1410 31300 1478 31356
rect 1534 31300 1602 31356
rect 1658 31300 1726 31356
rect 1782 31300 1850 31356
rect 1906 31300 2000 31356
rect 0 31232 2000 31300
rect 0 31176 114 31232
rect 170 31176 238 31232
rect 294 31176 362 31232
rect 418 31176 486 31232
rect 542 31176 610 31232
rect 666 31176 734 31232
rect 790 31176 858 31232
rect 914 31176 982 31232
rect 1038 31176 1106 31232
rect 1162 31176 1230 31232
rect 1286 31176 1354 31232
rect 1410 31176 1478 31232
rect 1534 31176 1602 31232
rect 1658 31176 1726 31232
rect 1782 31176 1850 31232
rect 1906 31176 2000 31232
rect 0 31108 2000 31176
rect 0 31052 114 31108
rect 170 31052 238 31108
rect 294 31052 362 31108
rect 418 31052 486 31108
rect 542 31052 610 31108
rect 666 31052 734 31108
rect 790 31052 858 31108
rect 914 31052 982 31108
rect 1038 31052 1106 31108
rect 1162 31052 1230 31108
rect 1286 31052 1354 31108
rect 1410 31052 1478 31108
rect 1534 31052 1602 31108
rect 1658 31052 1726 31108
rect 1782 31052 1850 31108
rect 1906 31052 2000 31108
rect 0 30984 2000 31052
rect 0 30928 114 30984
rect 170 30928 238 30984
rect 294 30928 362 30984
rect 418 30928 486 30984
rect 542 30928 610 30984
rect 666 30928 734 30984
rect 790 30928 858 30984
rect 914 30928 982 30984
rect 1038 30928 1106 30984
rect 1162 30928 1230 30984
rect 1286 30928 1354 30984
rect 1410 30928 1478 30984
rect 1534 30928 1602 30984
rect 1658 30928 1726 30984
rect 1782 30928 1850 30984
rect 1906 30928 2000 30984
rect 0 30860 2000 30928
rect 0 30804 114 30860
rect 170 30804 238 30860
rect 294 30804 362 30860
rect 418 30804 486 30860
rect 542 30804 610 30860
rect 666 30804 734 30860
rect 790 30804 858 30860
rect 914 30804 982 30860
rect 1038 30804 1106 30860
rect 1162 30804 1230 30860
rect 1286 30804 1354 30860
rect 1410 30804 1478 30860
rect 1534 30804 1602 30860
rect 1658 30804 1726 30860
rect 1782 30804 1850 30860
rect 1906 30804 2000 30860
rect 0 30736 2000 30804
rect 0 30680 114 30736
rect 170 30680 238 30736
rect 294 30680 362 30736
rect 418 30680 486 30736
rect 542 30680 610 30736
rect 666 30680 734 30736
rect 790 30680 858 30736
rect 914 30680 982 30736
rect 1038 30680 1106 30736
rect 1162 30680 1230 30736
rect 1286 30680 1354 30736
rect 1410 30680 1478 30736
rect 1534 30680 1602 30736
rect 1658 30680 1726 30736
rect 1782 30680 1850 30736
rect 1906 30680 2000 30736
rect 0 30612 2000 30680
rect 0 30556 114 30612
rect 170 30556 238 30612
rect 294 30556 362 30612
rect 418 30556 486 30612
rect 542 30556 610 30612
rect 666 30556 734 30612
rect 790 30556 858 30612
rect 914 30556 982 30612
rect 1038 30556 1106 30612
rect 1162 30556 1230 30612
rect 1286 30556 1354 30612
rect 1410 30556 1478 30612
rect 1534 30556 1602 30612
rect 1658 30556 1726 30612
rect 1782 30556 1850 30612
rect 1906 30556 2000 30612
rect 0 30488 2000 30556
rect 0 30432 114 30488
rect 170 30432 238 30488
rect 294 30432 362 30488
rect 418 30432 486 30488
rect 542 30432 610 30488
rect 666 30432 734 30488
rect 790 30432 858 30488
rect 914 30432 982 30488
rect 1038 30432 1106 30488
rect 1162 30432 1230 30488
rect 1286 30432 1354 30488
rect 1410 30432 1478 30488
rect 1534 30432 1602 30488
rect 1658 30432 1726 30488
rect 1782 30432 1850 30488
rect 1906 30432 2000 30488
rect 0 30364 2000 30432
rect 0 30308 114 30364
rect 170 30308 238 30364
rect 294 30308 362 30364
rect 418 30308 486 30364
rect 542 30308 610 30364
rect 666 30308 734 30364
rect 790 30308 858 30364
rect 914 30308 982 30364
rect 1038 30308 1106 30364
rect 1162 30308 1230 30364
rect 1286 30308 1354 30364
rect 1410 30308 1478 30364
rect 1534 30308 1602 30364
rect 1658 30308 1726 30364
rect 1782 30308 1850 30364
rect 1906 30308 2000 30364
rect 0 30240 2000 30308
rect 0 30184 114 30240
rect 170 30184 238 30240
rect 294 30184 362 30240
rect 418 30184 486 30240
rect 542 30184 610 30240
rect 666 30184 734 30240
rect 790 30184 858 30240
rect 914 30184 982 30240
rect 1038 30184 1106 30240
rect 1162 30184 1230 30240
rect 1286 30184 1354 30240
rect 1410 30184 1478 30240
rect 1534 30184 1602 30240
rect 1658 30184 1726 30240
rect 1782 30184 1850 30240
rect 1906 30184 2000 30240
rect 0 30000 2000 30184
rect 0 29643 2000 29800
rect 0 29587 114 29643
rect 170 29587 238 29643
rect 294 29587 362 29643
rect 418 29587 486 29643
rect 542 29587 610 29643
rect 666 29587 734 29643
rect 790 29587 858 29643
rect 914 29587 982 29643
rect 1038 29587 1106 29643
rect 1162 29587 1230 29643
rect 1286 29587 1354 29643
rect 1410 29587 1478 29643
rect 1534 29587 1602 29643
rect 1658 29587 1726 29643
rect 1782 29587 1850 29643
rect 1906 29587 2000 29643
rect 0 29519 2000 29587
rect 0 29463 114 29519
rect 170 29463 238 29519
rect 294 29463 362 29519
rect 418 29463 486 29519
rect 542 29463 610 29519
rect 666 29463 734 29519
rect 790 29463 858 29519
rect 914 29463 982 29519
rect 1038 29463 1106 29519
rect 1162 29463 1230 29519
rect 1286 29463 1354 29519
rect 1410 29463 1478 29519
rect 1534 29463 1602 29519
rect 1658 29463 1726 29519
rect 1782 29463 1850 29519
rect 1906 29463 2000 29519
rect 0 29395 2000 29463
rect 0 29339 114 29395
rect 170 29339 238 29395
rect 294 29339 362 29395
rect 418 29339 486 29395
rect 542 29339 610 29395
rect 666 29339 734 29395
rect 790 29339 858 29395
rect 914 29339 982 29395
rect 1038 29339 1106 29395
rect 1162 29339 1230 29395
rect 1286 29339 1354 29395
rect 1410 29339 1478 29395
rect 1534 29339 1602 29395
rect 1658 29339 1726 29395
rect 1782 29339 1850 29395
rect 1906 29339 2000 29395
rect 0 29271 2000 29339
rect 0 29215 114 29271
rect 170 29215 238 29271
rect 294 29215 362 29271
rect 418 29215 486 29271
rect 542 29215 610 29271
rect 666 29215 734 29271
rect 790 29215 858 29271
rect 914 29215 982 29271
rect 1038 29215 1106 29271
rect 1162 29215 1230 29271
rect 1286 29215 1354 29271
rect 1410 29215 1478 29271
rect 1534 29215 1602 29271
rect 1658 29215 1726 29271
rect 1782 29215 1850 29271
rect 1906 29215 2000 29271
rect 0 29147 2000 29215
rect 0 29091 114 29147
rect 170 29091 238 29147
rect 294 29091 362 29147
rect 418 29091 486 29147
rect 542 29091 610 29147
rect 666 29091 734 29147
rect 790 29091 858 29147
rect 914 29091 982 29147
rect 1038 29091 1106 29147
rect 1162 29091 1230 29147
rect 1286 29091 1354 29147
rect 1410 29091 1478 29147
rect 1534 29091 1602 29147
rect 1658 29091 1726 29147
rect 1782 29091 1850 29147
rect 1906 29091 2000 29147
rect 0 29023 2000 29091
rect 0 28967 114 29023
rect 170 28967 238 29023
rect 294 28967 362 29023
rect 418 28967 486 29023
rect 542 28967 610 29023
rect 666 28967 734 29023
rect 790 28967 858 29023
rect 914 28967 982 29023
rect 1038 28967 1106 29023
rect 1162 28967 1230 29023
rect 1286 28967 1354 29023
rect 1410 28967 1478 29023
rect 1534 28967 1602 29023
rect 1658 28967 1726 29023
rect 1782 28967 1850 29023
rect 1906 28967 2000 29023
rect 0 28899 2000 28967
rect 0 28843 114 28899
rect 170 28843 238 28899
rect 294 28843 362 28899
rect 418 28843 486 28899
rect 542 28843 610 28899
rect 666 28843 734 28899
rect 790 28843 858 28899
rect 914 28843 982 28899
rect 1038 28843 1106 28899
rect 1162 28843 1230 28899
rect 1286 28843 1354 28899
rect 1410 28843 1478 28899
rect 1534 28843 1602 28899
rect 1658 28843 1726 28899
rect 1782 28843 1850 28899
rect 1906 28843 2000 28899
rect 0 28775 2000 28843
rect 0 28719 114 28775
rect 170 28719 238 28775
rect 294 28719 362 28775
rect 418 28719 486 28775
rect 542 28719 610 28775
rect 666 28719 734 28775
rect 790 28719 858 28775
rect 914 28719 982 28775
rect 1038 28719 1106 28775
rect 1162 28719 1230 28775
rect 1286 28719 1354 28775
rect 1410 28719 1478 28775
rect 1534 28719 1602 28775
rect 1658 28719 1726 28775
rect 1782 28719 1850 28775
rect 1906 28719 2000 28775
rect 0 28651 2000 28719
rect 0 28595 114 28651
rect 170 28595 238 28651
rect 294 28595 362 28651
rect 418 28595 486 28651
rect 542 28595 610 28651
rect 666 28595 734 28651
rect 790 28595 858 28651
rect 914 28595 982 28651
rect 1038 28595 1106 28651
rect 1162 28595 1230 28651
rect 1286 28595 1354 28651
rect 1410 28595 1478 28651
rect 1534 28595 1602 28651
rect 1658 28595 1726 28651
rect 1782 28595 1850 28651
rect 1906 28595 2000 28651
rect 0 28527 2000 28595
rect 0 28471 114 28527
rect 170 28471 238 28527
rect 294 28471 362 28527
rect 418 28471 486 28527
rect 542 28471 610 28527
rect 666 28471 734 28527
rect 790 28471 858 28527
rect 914 28471 982 28527
rect 1038 28471 1106 28527
rect 1162 28471 1230 28527
rect 1286 28471 1354 28527
rect 1410 28471 1478 28527
rect 1534 28471 1602 28527
rect 1658 28471 1726 28527
rect 1782 28471 1850 28527
rect 1906 28471 2000 28527
rect 0 28403 2000 28471
rect 0 28347 114 28403
rect 170 28347 238 28403
rect 294 28347 362 28403
rect 418 28347 486 28403
rect 542 28347 610 28403
rect 666 28347 734 28403
rect 790 28347 858 28403
rect 914 28347 982 28403
rect 1038 28347 1106 28403
rect 1162 28347 1230 28403
rect 1286 28347 1354 28403
rect 1410 28347 1478 28403
rect 1534 28347 1602 28403
rect 1658 28347 1726 28403
rect 1782 28347 1850 28403
rect 1906 28347 2000 28403
rect 0 28279 2000 28347
rect 0 28223 114 28279
rect 170 28223 238 28279
rect 294 28223 362 28279
rect 418 28223 486 28279
rect 542 28223 610 28279
rect 666 28223 734 28279
rect 790 28223 858 28279
rect 914 28223 982 28279
rect 1038 28223 1106 28279
rect 1162 28223 1230 28279
rect 1286 28223 1354 28279
rect 1410 28223 1478 28279
rect 1534 28223 1602 28279
rect 1658 28223 1726 28279
rect 1782 28223 1850 28279
rect 1906 28223 2000 28279
rect 0 28155 2000 28223
rect 0 28099 114 28155
rect 170 28099 238 28155
rect 294 28099 362 28155
rect 418 28099 486 28155
rect 542 28099 610 28155
rect 666 28099 734 28155
rect 790 28099 858 28155
rect 914 28099 982 28155
rect 1038 28099 1106 28155
rect 1162 28099 1230 28155
rect 1286 28099 1354 28155
rect 1410 28099 1478 28155
rect 1534 28099 1602 28155
rect 1658 28099 1726 28155
rect 1782 28099 1850 28155
rect 1906 28099 2000 28155
rect 0 28031 2000 28099
rect 0 27975 114 28031
rect 170 27975 238 28031
rect 294 27975 362 28031
rect 418 27975 486 28031
rect 542 27975 610 28031
rect 666 27975 734 28031
rect 790 27975 858 28031
rect 914 27975 982 28031
rect 1038 27975 1106 28031
rect 1162 27975 1230 28031
rect 1286 27975 1354 28031
rect 1410 27975 1478 28031
rect 1534 27975 1602 28031
rect 1658 27975 1726 28031
rect 1782 27975 1850 28031
rect 1906 27975 2000 28031
rect 0 27907 2000 27975
rect 0 27851 114 27907
rect 170 27851 238 27907
rect 294 27851 362 27907
rect 418 27851 486 27907
rect 542 27851 610 27907
rect 666 27851 734 27907
rect 790 27851 858 27907
rect 914 27851 982 27907
rect 1038 27851 1106 27907
rect 1162 27851 1230 27907
rect 1286 27851 1354 27907
rect 1410 27851 1478 27907
rect 1534 27851 1602 27907
rect 1658 27851 1726 27907
rect 1782 27851 1850 27907
rect 1906 27851 2000 27907
rect 0 27783 2000 27851
rect 0 27727 114 27783
rect 170 27727 238 27783
rect 294 27727 362 27783
rect 418 27727 486 27783
rect 542 27727 610 27783
rect 666 27727 734 27783
rect 790 27727 858 27783
rect 914 27727 982 27783
rect 1038 27727 1106 27783
rect 1162 27727 1230 27783
rect 1286 27727 1354 27783
rect 1410 27727 1478 27783
rect 1534 27727 1602 27783
rect 1658 27727 1726 27783
rect 1782 27727 1850 27783
rect 1906 27727 2000 27783
rect 0 27659 2000 27727
rect 0 27603 114 27659
rect 170 27603 238 27659
rect 294 27603 362 27659
rect 418 27603 486 27659
rect 542 27603 610 27659
rect 666 27603 734 27659
rect 790 27603 858 27659
rect 914 27603 982 27659
rect 1038 27603 1106 27659
rect 1162 27603 1230 27659
rect 1286 27603 1354 27659
rect 1410 27603 1478 27659
rect 1534 27603 1602 27659
rect 1658 27603 1726 27659
rect 1782 27603 1850 27659
rect 1906 27603 2000 27659
rect 0 27535 2000 27603
rect 0 27479 114 27535
rect 170 27479 238 27535
rect 294 27479 362 27535
rect 418 27479 486 27535
rect 542 27479 610 27535
rect 666 27479 734 27535
rect 790 27479 858 27535
rect 914 27479 982 27535
rect 1038 27479 1106 27535
rect 1162 27479 1230 27535
rect 1286 27479 1354 27535
rect 1410 27479 1478 27535
rect 1534 27479 1602 27535
rect 1658 27479 1726 27535
rect 1782 27479 1850 27535
rect 1906 27479 2000 27535
rect 0 27411 2000 27479
rect 0 27355 114 27411
rect 170 27355 238 27411
rect 294 27355 362 27411
rect 418 27355 486 27411
rect 542 27355 610 27411
rect 666 27355 734 27411
rect 790 27355 858 27411
rect 914 27355 982 27411
rect 1038 27355 1106 27411
rect 1162 27355 1230 27411
rect 1286 27355 1354 27411
rect 1410 27355 1478 27411
rect 1534 27355 1602 27411
rect 1658 27355 1726 27411
rect 1782 27355 1850 27411
rect 1906 27355 2000 27411
rect 0 27287 2000 27355
rect 0 27231 114 27287
rect 170 27231 238 27287
rect 294 27231 362 27287
rect 418 27231 486 27287
rect 542 27231 610 27287
rect 666 27231 734 27287
rect 790 27231 858 27287
rect 914 27231 982 27287
rect 1038 27231 1106 27287
rect 1162 27231 1230 27287
rect 1286 27231 1354 27287
rect 1410 27231 1478 27287
rect 1534 27231 1602 27287
rect 1658 27231 1726 27287
rect 1782 27231 1850 27287
rect 1906 27231 2000 27287
rect 0 27163 2000 27231
rect 0 27107 114 27163
rect 170 27107 238 27163
rect 294 27107 362 27163
rect 418 27107 486 27163
rect 542 27107 610 27163
rect 666 27107 734 27163
rect 790 27107 858 27163
rect 914 27107 982 27163
rect 1038 27107 1106 27163
rect 1162 27107 1230 27163
rect 1286 27107 1354 27163
rect 1410 27107 1478 27163
rect 1534 27107 1602 27163
rect 1658 27107 1726 27163
rect 1782 27107 1850 27163
rect 1906 27107 2000 27163
rect 0 27039 2000 27107
rect 0 26983 114 27039
rect 170 26983 238 27039
rect 294 26983 362 27039
rect 418 26983 486 27039
rect 542 26983 610 27039
rect 666 26983 734 27039
rect 790 26983 858 27039
rect 914 26983 982 27039
rect 1038 26983 1106 27039
rect 1162 26983 1230 27039
rect 1286 26983 1354 27039
rect 1410 26983 1478 27039
rect 1534 26983 1602 27039
rect 1658 26983 1726 27039
rect 1782 26983 1850 27039
rect 1906 26983 2000 27039
rect 0 26800 2000 26983
rect 0 26501 2000 26600
rect 0 26445 114 26501
rect 170 26445 238 26501
rect 294 26445 362 26501
rect 418 26445 486 26501
rect 542 26445 610 26501
rect 666 26445 734 26501
rect 790 26445 858 26501
rect 914 26445 982 26501
rect 1038 26445 1106 26501
rect 1162 26445 1230 26501
rect 1286 26445 1354 26501
rect 1410 26445 1478 26501
rect 1534 26445 1602 26501
rect 1658 26445 1726 26501
rect 1782 26445 1850 26501
rect 1906 26445 2000 26501
rect 0 26377 2000 26445
rect 0 26321 114 26377
rect 170 26321 238 26377
rect 294 26321 362 26377
rect 418 26321 486 26377
rect 542 26321 610 26377
rect 666 26321 734 26377
rect 790 26321 858 26377
rect 914 26321 982 26377
rect 1038 26321 1106 26377
rect 1162 26321 1230 26377
rect 1286 26321 1354 26377
rect 1410 26321 1478 26377
rect 1534 26321 1602 26377
rect 1658 26321 1726 26377
rect 1782 26321 1850 26377
rect 1906 26321 2000 26377
rect 0 26253 2000 26321
rect 0 26197 114 26253
rect 170 26197 238 26253
rect 294 26197 362 26253
rect 418 26197 486 26253
rect 542 26197 610 26253
rect 666 26197 734 26253
rect 790 26197 858 26253
rect 914 26197 982 26253
rect 1038 26197 1106 26253
rect 1162 26197 1230 26253
rect 1286 26197 1354 26253
rect 1410 26197 1478 26253
rect 1534 26197 1602 26253
rect 1658 26197 1726 26253
rect 1782 26197 1850 26253
rect 1906 26197 2000 26253
rect 0 26129 2000 26197
rect 0 26073 114 26129
rect 170 26073 238 26129
rect 294 26073 362 26129
rect 418 26073 486 26129
rect 542 26073 610 26129
rect 666 26073 734 26129
rect 790 26073 858 26129
rect 914 26073 982 26129
rect 1038 26073 1106 26129
rect 1162 26073 1230 26129
rect 1286 26073 1354 26129
rect 1410 26073 1478 26129
rect 1534 26073 1602 26129
rect 1658 26073 1726 26129
rect 1782 26073 1850 26129
rect 1906 26073 2000 26129
rect 0 26005 2000 26073
rect 0 25949 114 26005
rect 170 25949 238 26005
rect 294 25949 362 26005
rect 418 25949 486 26005
rect 542 25949 610 26005
rect 666 25949 734 26005
rect 790 25949 858 26005
rect 914 25949 982 26005
rect 1038 25949 1106 26005
rect 1162 25949 1230 26005
rect 1286 25949 1354 26005
rect 1410 25949 1478 26005
rect 1534 25949 1602 26005
rect 1658 25949 1726 26005
rect 1782 25949 1850 26005
rect 1906 25949 2000 26005
rect 0 25881 2000 25949
rect 0 25825 114 25881
rect 170 25825 238 25881
rect 294 25825 362 25881
rect 418 25825 486 25881
rect 542 25825 610 25881
rect 666 25825 734 25881
rect 790 25825 858 25881
rect 914 25825 982 25881
rect 1038 25825 1106 25881
rect 1162 25825 1230 25881
rect 1286 25825 1354 25881
rect 1410 25825 1478 25881
rect 1534 25825 1602 25881
rect 1658 25825 1726 25881
rect 1782 25825 1850 25881
rect 1906 25825 2000 25881
rect 0 25757 2000 25825
rect 0 25701 114 25757
rect 170 25701 238 25757
rect 294 25701 362 25757
rect 418 25701 486 25757
rect 542 25701 610 25757
rect 666 25701 734 25757
rect 790 25701 858 25757
rect 914 25701 982 25757
rect 1038 25701 1106 25757
rect 1162 25701 1230 25757
rect 1286 25701 1354 25757
rect 1410 25701 1478 25757
rect 1534 25701 1602 25757
rect 1658 25701 1726 25757
rect 1782 25701 1850 25757
rect 1906 25701 2000 25757
rect 0 25633 2000 25701
rect 0 25577 114 25633
rect 170 25577 238 25633
rect 294 25577 362 25633
rect 418 25577 486 25633
rect 542 25577 610 25633
rect 666 25577 734 25633
rect 790 25577 858 25633
rect 914 25577 982 25633
rect 1038 25577 1106 25633
rect 1162 25577 1230 25633
rect 1286 25577 1354 25633
rect 1410 25577 1478 25633
rect 1534 25577 1602 25633
rect 1658 25577 1726 25633
rect 1782 25577 1850 25633
rect 1906 25577 2000 25633
rect 0 25509 2000 25577
rect 0 25453 114 25509
rect 170 25453 238 25509
rect 294 25453 362 25509
rect 418 25453 486 25509
rect 542 25453 610 25509
rect 666 25453 734 25509
rect 790 25453 858 25509
rect 914 25453 982 25509
rect 1038 25453 1106 25509
rect 1162 25453 1230 25509
rect 1286 25453 1354 25509
rect 1410 25453 1478 25509
rect 1534 25453 1602 25509
rect 1658 25453 1726 25509
rect 1782 25453 1850 25509
rect 1906 25453 2000 25509
rect 0 25385 2000 25453
rect 0 25329 114 25385
rect 170 25329 238 25385
rect 294 25329 362 25385
rect 418 25329 486 25385
rect 542 25329 610 25385
rect 666 25329 734 25385
rect 790 25329 858 25385
rect 914 25329 982 25385
rect 1038 25329 1106 25385
rect 1162 25329 1230 25385
rect 1286 25329 1354 25385
rect 1410 25329 1478 25385
rect 1534 25329 1602 25385
rect 1658 25329 1726 25385
rect 1782 25329 1850 25385
rect 1906 25329 2000 25385
rect 0 25200 2000 25329
rect 0 24888 2000 25000
rect 0 24832 114 24888
rect 170 24832 238 24888
rect 294 24832 362 24888
rect 418 24832 486 24888
rect 542 24832 610 24888
rect 666 24832 734 24888
rect 790 24832 858 24888
rect 914 24832 982 24888
rect 1038 24832 1106 24888
rect 1162 24832 1230 24888
rect 1286 24832 1354 24888
rect 1410 24832 1478 24888
rect 1534 24832 1602 24888
rect 1658 24832 1726 24888
rect 1782 24832 1850 24888
rect 1906 24832 2000 24888
rect 0 24764 2000 24832
rect 0 24708 114 24764
rect 170 24708 238 24764
rect 294 24708 362 24764
rect 418 24708 486 24764
rect 542 24708 610 24764
rect 666 24708 734 24764
rect 790 24708 858 24764
rect 914 24708 982 24764
rect 1038 24708 1106 24764
rect 1162 24708 1230 24764
rect 1286 24708 1354 24764
rect 1410 24708 1478 24764
rect 1534 24708 1602 24764
rect 1658 24708 1726 24764
rect 1782 24708 1850 24764
rect 1906 24708 2000 24764
rect 0 24640 2000 24708
rect 0 24584 114 24640
rect 170 24584 238 24640
rect 294 24584 362 24640
rect 418 24584 486 24640
rect 542 24584 610 24640
rect 666 24584 734 24640
rect 790 24584 858 24640
rect 914 24584 982 24640
rect 1038 24584 1106 24640
rect 1162 24584 1230 24640
rect 1286 24584 1354 24640
rect 1410 24584 1478 24640
rect 1534 24584 1602 24640
rect 1658 24584 1726 24640
rect 1782 24584 1850 24640
rect 1906 24584 2000 24640
rect 0 24516 2000 24584
rect 0 24460 114 24516
rect 170 24460 238 24516
rect 294 24460 362 24516
rect 418 24460 486 24516
rect 542 24460 610 24516
rect 666 24460 734 24516
rect 790 24460 858 24516
rect 914 24460 982 24516
rect 1038 24460 1106 24516
rect 1162 24460 1230 24516
rect 1286 24460 1354 24516
rect 1410 24460 1478 24516
rect 1534 24460 1602 24516
rect 1658 24460 1726 24516
rect 1782 24460 1850 24516
rect 1906 24460 2000 24516
rect 0 24392 2000 24460
rect 0 24336 114 24392
rect 170 24336 238 24392
rect 294 24336 362 24392
rect 418 24336 486 24392
rect 542 24336 610 24392
rect 666 24336 734 24392
rect 790 24336 858 24392
rect 914 24336 982 24392
rect 1038 24336 1106 24392
rect 1162 24336 1230 24392
rect 1286 24336 1354 24392
rect 1410 24336 1478 24392
rect 1534 24336 1602 24392
rect 1658 24336 1726 24392
rect 1782 24336 1850 24392
rect 1906 24336 2000 24392
rect 0 24268 2000 24336
rect 0 24212 114 24268
rect 170 24212 238 24268
rect 294 24212 362 24268
rect 418 24212 486 24268
rect 542 24212 610 24268
rect 666 24212 734 24268
rect 790 24212 858 24268
rect 914 24212 982 24268
rect 1038 24212 1106 24268
rect 1162 24212 1230 24268
rect 1286 24212 1354 24268
rect 1410 24212 1478 24268
rect 1534 24212 1602 24268
rect 1658 24212 1726 24268
rect 1782 24212 1850 24268
rect 1906 24212 2000 24268
rect 0 24144 2000 24212
rect 0 24088 114 24144
rect 170 24088 238 24144
rect 294 24088 362 24144
rect 418 24088 486 24144
rect 542 24088 610 24144
rect 666 24088 734 24144
rect 790 24088 858 24144
rect 914 24088 982 24144
rect 1038 24088 1106 24144
rect 1162 24088 1230 24144
rect 1286 24088 1354 24144
rect 1410 24088 1478 24144
rect 1534 24088 1602 24144
rect 1658 24088 1726 24144
rect 1782 24088 1850 24144
rect 1906 24088 2000 24144
rect 0 24020 2000 24088
rect 0 23964 114 24020
rect 170 23964 238 24020
rect 294 23964 362 24020
rect 418 23964 486 24020
rect 542 23964 610 24020
rect 666 23964 734 24020
rect 790 23964 858 24020
rect 914 23964 982 24020
rect 1038 23964 1106 24020
rect 1162 23964 1230 24020
rect 1286 23964 1354 24020
rect 1410 23964 1478 24020
rect 1534 23964 1602 24020
rect 1658 23964 1726 24020
rect 1782 23964 1850 24020
rect 1906 23964 2000 24020
rect 0 23896 2000 23964
rect 0 23840 114 23896
rect 170 23840 238 23896
rect 294 23840 362 23896
rect 418 23840 486 23896
rect 542 23840 610 23896
rect 666 23840 734 23896
rect 790 23840 858 23896
rect 914 23840 982 23896
rect 1038 23840 1106 23896
rect 1162 23840 1230 23896
rect 1286 23840 1354 23896
rect 1410 23840 1478 23896
rect 1534 23840 1602 23896
rect 1658 23840 1726 23896
rect 1782 23840 1850 23896
rect 1906 23840 2000 23896
rect 0 23772 2000 23840
rect 0 23716 114 23772
rect 170 23716 238 23772
rect 294 23716 362 23772
rect 418 23716 486 23772
rect 542 23716 610 23772
rect 666 23716 734 23772
rect 790 23716 858 23772
rect 914 23716 982 23772
rect 1038 23716 1106 23772
rect 1162 23716 1230 23772
rect 1286 23716 1354 23772
rect 1410 23716 1478 23772
rect 1534 23716 1602 23772
rect 1658 23716 1726 23772
rect 1782 23716 1850 23772
rect 1906 23716 2000 23772
rect 0 23600 2000 23716
rect 0 23234 2000 23400
rect 0 23178 114 23234
rect 170 23178 238 23234
rect 294 23178 362 23234
rect 418 23178 486 23234
rect 542 23178 610 23234
rect 666 23178 734 23234
rect 790 23178 858 23234
rect 914 23178 982 23234
rect 1038 23178 1106 23234
rect 1162 23178 1230 23234
rect 1286 23178 1354 23234
rect 1410 23178 1478 23234
rect 1534 23178 1602 23234
rect 1658 23178 1726 23234
rect 1782 23178 1850 23234
rect 1906 23178 2000 23234
rect 0 23110 2000 23178
rect 0 23054 114 23110
rect 170 23054 238 23110
rect 294 23054 362 23110
rect 418 23054 486 23110
rect 542 23054 610 23110
rect 666 23054 734 23110
rect 790 23054 858 23110
rect 914 23054 982 23110
rect 1038 23054 1106 23110
rect 1162 23054 1230 23110
rect 1286 23054 1354 23110
rect 1410 23054 1478 23110
rect 1534 23054 1602 23110
rect 1658 23054 1726 23110
rect 1782 23054 1850 23110
rect 1906 23054 2000 23110
rect 0 22986 2000 23054
rect 0 22930 114 22986
rect 170 22930 238 22986
rect 294 22930 362 22986
rect 418 22930 486 22986
rect 542 22930 610 22986
rect 666 22930 734 22986
rect 790 22930 858 22986
rect 914 22930 982 22986
rect 1038 22930 1106 22986
rect 1162 22930 1230 22986
rect 1286 22930 1354 22986
rect 1410 22930 1478 22986
rect 1534 22930 1602 22986
rect 1658 22930 1726 22986
rect 1782 22930 1850 22986
rect 1906 22930 2000 22986
rect 0 22862 2000 22930
rect 0 22806 114 22862
rect 170 22806 238 22862
rect 294 22806 362 22862
rect 418 22806 486 22862
rect 542 22806 610 22862
rect 666 22806 734 22862
rect 790 22806 858 22862
rect 914 22806 982 22862
rect 1038 22806 1106 22862
rect 1162 22806 1230 22862
rect 1286 22806 1354 22862
rect 1410 22806 1478 22862
rect 1534 22806 1602 22862
rect 1658 22806 1726 22862
rect 1782 22806 1850 22862
rect 1906 22806 2000 22862
rect 0 22738 2000 22806
rect 0 22682 114 22738
rect 170 22682 238 22738
rect 294 22682 362 22738
rect 418 22682 486 22738
rect 542 22682 610 22738
rect 666 22682 734 22738
rect 790 22682 858 22738
rect 914 22682 982 22738
rect 1038 22682 1106 22738
rect 1162 22682 1230 22738
rect 1286 22682 1354 22738
rect 1410 22682 1478 22738
rect 1534 22682 1602 22738
rect 1658 22682 1726 22738
rect 1782 22682 1850 22738
rect 1906 22682 2000 22738
rect 0 22614 2000 22682
rect 0 22558 114 22614
rect 170 22558 238 22614
rect 294 22558 362 22614
rect 418 22558 486 22614
rect 542 22558 610 22614
rect 666 22558 734 22614
rect 790 22558 858 22614
rect 914 22558 982 22614
rect 1038 22558 1106 22614
rect 1162 22558 1230 22614
rect 1286 22558 1354 22614
rect 1410 22558 1478 22614
rect 1534 22558 1602 22614
rect 1658 22558 1726 22614
rect 1782 22558 1850 22614
rect 1906 22558 2000 22614
rect 0 22490 2000 22558
rect 0 22434 114 22490
rect 170 22434 238 22490
rect 294 22434 362 22490
rect 418 22434 486 22490
rect 542 22434 610 22490
rect 666 22434 734 22490
rect 790 22434 858 22490
rect 914 22434 982 22490
rect 1038 22434 1106 22490
rect 1162 22434 1230 22490
rect 1286 22434 1354 22490
rect 1410 22434 1478 22490
rect 1534 22434 1602 22490
rect 1658 22434 1726 22490
rect 1782 22434 1850 22490
rect 1906 22434 2000 22490
rect 0 22366 2000 22434
rect 0 22310 114 22366
rect 170 22310 238 22366
rect 294 22310 362 22366
rect 418 22310 486 22366
rect 542 22310 610 22366
rect 666 22310 734 22366
rect 790 22310 858 22366
rect 914 22310 982 22366
rect 1038 22310 1106 22366
rect 1162 22310 1230 22366
rect 1286 22310 1354 22366
rect 1410 22310 1478 22366
rect 1534 22310 1602 22366
rect 1658 22310 1726 22366
rect 1782 22310 1850 22366
rect 1906 22310 2000 22366
rect 0 22242 2000 22310
rect 0 22186 114 22242
rect 170 22186 238 22242
rect 294 22186 362 22242
rect 418 22186 486 22242
rect 542 22186 610 22242
rect 666 22186 734 22242
rect 790 22186 858 22242
rect 914 22186 982 22242
rect 1038 22186 1106 22242
rect 1162 22186 1230 22242
rect 1286 22186 1354 22242
rect 1410 22186 1478 22242
rect 1534 22186 1602 22242
rect 1658 22186 1726 22242
rect 1782 22186 1850 22242
rect 1906 22186 2000 22242
rect 0 22118 2000 22186
rect 0 22062 114 22118
rect 170 22062 238 22118
rect 294 22062 362 22118
rect 418 22062 486 22118
rect 542 22062 610 22118
rect 666 22062 734 22118
rect 790 22062 858 22118
rect 914 22062 982 22118
rect 1038 22062 1106 22118
rect 1162 22062 1230 22118
rect 1286 22062 1354 22118
rect 1410 22062 1478 22118
rect 1534 22062 1602 22118
rect 1658 22062 1726 22118
rect 1782 22062 1850 22118
rect 1906 22062 2000 22118
rect 0 21994 2000 22062
rect 0 21938 114 21994
rect 170 21938 238 21994
rect 294 21938 362 21994
rect 418 21938 486 21994
rect 542 21938 610 21994
rect 666 21938 734 21994
rect 790 21938 858 21994
rect 914 21938 982 21994
rect 1038 21938 1106 21994
rect 1162 21938 1230 21994
rect 1286 21938 1354 21994
rect 1410 21938 1478 21994
rect 1534 21938 1602 21994
rect 1658 21938 1726 21994
rect 1782 21938 1850 21994
rect 1906 21938 2000 21994
rect 0 21870 2000 21938
rect 0 21814 114 21870
rect 170 21814 238 21870
rect 294 21814 362 21870
rect 418 21814 486 21870
rect 542 21814 610 21870
rect 666 21814 734 21870
rect 790 21814 858 21870
rect 914 21814 982 21870
rect 1038 21814 1106 21870
rect 1162 21814 1230 21870
rect 1286 21814 1354 21870
rect 1410 21814 1478 21870
rect 1534 21814 1602 21870
rect 1658 21814 1726 21870
rect 1782 21814 1850 21870
rect 1906 21814 2000 21870
rect 0 21746 2000 21814
rect 0 21690 114 21746
rect 170 21690 238 21746
rect 294 21690 362 21746
rect 418 21690 486 21746
rect 542 21690 610 21746
rect 666 21690 734 21746
rect 790 21690 858 21746
rect 914 21690 982 21746
rect 1038 21690 1106 21746
rect 1162 21690 1230 21746
rect 1286 21690 1354 21746
rect 1410 21690 1478 21746
rect 1534 21690 1602 21746
rect 1658 21690 1726 21746
rect 1782 21690 1850 21746
rect 1906 21690 2000 21746
rect 0 21622 2000 21690
rect 0 21566 114 21622
rect 170 21566 238 21622
rect 294 21566 362 21622
rect 418 21566 486 21622
rect 542 21566 610 21622
rect 666 21566 734 21622
rect 790 21566 858 21622
rect 914 21566 982 21622
rect 1038 21566 1106 21622
rect 1162 21566 1230 21622
rect 1286 21566 1354 21622
rect 1410 21566 1478 21622
rect 1534 21566 1602 21622
rect 1658 21566 1726 21622
rect 1782 21566 1850 21622
rect 1906 21566 2000 21622
rect 0 21498 2000 21566
rect 0 21442 114 21498
rect 170 21442 238 21498
rect 294 21442 362 21498
rect 418 21442 486 21498
rect 542 21442 610 21498
rect 666 21442 734 21498
rect 790 21442 858 21498
rect 914 21442 982 21498
rect 1038 21442 1106 21498
rect 1162 21442 1230 21498
rect 1286 21442 1354 21498
rect 1410 21442 1478 21498
rect 1534 21442 1602 21498
rect 1658 21442 1726 21498
rect 1782 21442 1850 21498
rect 1906 21442 2000 21498
rect 0 21374 2000 21442
rect 0 21318 114 21374
rect 170 21318 238 21374
rect 294 21318 362 21374
rect 418 21318 486 21374
rect 542 21318 610 21374
rect 666 21318 734 21374
rect 790 21318 858 21374
rect 914 21318 982 21374
rect 1038 21318 1106 21374
rect 1162 21318 1230 21374
rect 1286 21318 1354 21374
rect 1410 21318 1478 21374
rect 1534 21318 1602 21374
rect 1658 21318 1726 21374
rect 1782 21318 1850 21374
rect 1906 21318 2000 21374
rect 0 21250 2000 21318
rect 0 21194 114 21250
rect 170 21194 238 21250
rect 294 21194 362 21250
rect 418 21194 486 21250
rect 542 21194 610 21250
rect 666 21194 734 21250
rect 790 21194 858 21250
rect 914 21194 982 21250
rect 1038 21194 1106 21250
rect 1162 21194 1230 21250
rect 1286 21194 1354 21250
rect 1410 21194 1478 21250
rect 1534 21194 1602 21250
rect 1658 21194 1726 21250
rect 1782 21194 1850 21250
rect 1906 21194 2000 21250
rect 0 21126 2000 21194
rect 0 21070 114 21126
rect 170 21070 238 21126
rect 294 21070 362 21126
rect 418 21070 486 21126
rect 542 21070 610 21126
rect 666 21070 734 21126
rect 790 21070 858 21126
rect 914 21070 982 21126
rect 1038 21070 1106 21126
rect 1162 21070 1230 21126
rect 1286 21070 1354 21126
rect 1410 21070 1478 21126
rect 1534 21070 1602 21126
rect 1658 21070 1726 21126
rect 1782 21070 1850 21126
rect 1906 21070 2000 21126
rect 0 21002 2000 21070
rect 0 20946 114 21002
rect 170 20946 238 21002
rect 294 20946 362 21002
rect 418 20946 486 21002
rect 542 20946 610 21002
rect 666 20946 734 21002
rect 790 20946 858 21002
rect 914 20946 982 21002
rect 1038 20946 1106 21002
rect 1162 20946 1230 21002
rect 1286 20946 1354 21002
rect 1410 20946 1478 21002
rect 1534 20946 1602 21002
rect 1658 20946 1726 21002
rect 1782 20946 1850 21002
rect 1906 20946 2000 21002
rect 0 20878 2000 20946
rect 0 20822 114 20878
rect 170 20822 238 20878
rect 294 20822 362 20878
rect 418 20822 486 20878
rect 542 20822 610 20878
rect 666 20822 734 20878
rect 790 20822 858 20878
rect 914 20822 982 20878
rect 1038 20822 1106 20878
rect 1162 20822 1230 20878
rect 1286 20822 1354 20878
rect 1410 20822 1478 20878
rect 1534 20822 1602 20878
rect 1658 20822 1726 20878
rect 1782 20822 1850 20878
rect 1906 20822 2000 20878
rect 0 20754 2000 20822
rect 0 20698 114 20754
rect 170 20698 238 20754
rect 294 20698 362 20754
rect 418 20698 486 20754
rect 542 20698 610 20754
rect 666 20698 734 20754
rect 790 20698 858 20754
rect 914 20698 982 20754
rect 1038 20698 1106 20754
rect 1162 20698 1230 20754
rect 1286 20698 1354 20754
rect 1410 20698 1478 20754
rect 1534 20698 1602 20754
rect 1658 20698 1726 20754
rect 1782 20698 1850 20754
rect 1906 20698 2000 20754
rect 0 20630 2000 20698
rect 0 20574 114 20630
rect 170 20574 238 20630
rect 294 20574 362 20630
rect 418 20574 486 20630
rect 542 20574 610 20630
rect 666 20574 734 20630
rect 790 20574 858 20630
rect 914 20574 982 20630
rect 1038 20574 1106 20630
rect 1162 20574 1230 20630
rect 1286 20574 1354 20630
rect 1410 20574 1478 20630
rect 1534 20574 1602 20630
rect 1658 20574 1726 20630
rect 1782 20574 1850 20630
rect 1906 20574 2000 20630
rect 0 20400 2000 20574
rect 0 20023 2000 20200
rect 0 19967 114 20023
rect 170 19967 238 20023
rect 294 19967 362 20023
rect 418 19967 486 20023
rect 542 19967 610 20023
rect 666 19967 734 20023
rect 790 19967 858 20023
rect 914 19967 982 20023
rect 1038 19967 1106 20023
rect 1162 19967 1230 20023
rect 1286 19967 1354 20023
rect 1410 19967 1478 20023
rect 1534 19967 1602 20023
rect 1658 19967 1726 20023
rect 1782 19967 1850 20023
rect 1906 19967 2000 20023
rect 0 19899 2000 19967
rect 0 19843 114 19899
rect 170 19843 238 19899
rect 294 19843 362 19899
rect 418 19843 486 19899
rect 542 19843 610 19899
rect 666 19843 734 19899
rect 790 19843 858 19899
rect 914 19843 982 19899
rect 1038 19843 1106 19899
rect 1162 19843 1230 19899
rect 1286 19843 1354 19899
rect 1410 19843 1478 19899
rect 1534 19843 1602 19899
rect 1658 19843 1726 19899
rect 1782 19843 1850 19899
rect 1906 19843 2000 19899
rect 0 19775 2000 19843
rect 0 19719 114 19775
rect 170 19719 238 19775
rect 294 19719 362 19775
rect 418 19719 486 19775
rect 542 19719 610 19775
rect 666 19719 734 19775
rect 790 19719 858 19775
rect 914 19719 982 19775
rect 1038 19719 1106 19775
rect 1162 19719 1230 19775
rect 1286 19719 1354 19775
rect 1410 19719 1478 19775
rect 1534 19719 1602 19775
rect 1658 19719 1726 19775
rect 1782 19719 1850 19775
rect 1906 19719 2000 19775
rect 0 19651 2000 19719
rect 0 19595 114 19651
rect 170 19595 238 19651
rect 294 19595 362 19651
rect 418 19595 486 19651
rect 542 19595 610 19651
rect 666 19595 734 19651
rect 790 19595 858 19651
rect 914 19595 982 19651
rect 1038 19595 1106 19651
rect 1162 19595 1230 19651
rect 1286 19595 1354 19651
rect 1410 19595 1478 19651
rect 1534 19595 1602 19651
rect 1658 19595 1726 19651
rect 1782 19595 1850 19651
rect 1906 19595 2000 19651
rect 0 19527 2000 19595
rect 0 19471 114 19527
rect 170 19471 238 19527
rect 294 19471 362 19527
rect 418 19471 486 19527
rect 542 19471 610 19527
rect 666 19471 734 19527
rect 790 19471 858 19527
rect 914 19471 982 19527
rect 1038 19471 1106 19527
rect 1162 19471 1230 19527
rect 1286 19471 1354 19527
rect 1410 19471 1478 19527
rect 1534 19471 1602 19527
rect 1658 19471 1726 19527
rect 1782 19471 1850 19527
rect 1906 19471 2000 19527
rect 0 19403 2000 19471
rect 0 19347 114 19403
rect 170 19347 238 19403
rect 294 19347 362 19403
rect 418 19347 486 19403
rect 542 19347 610 19403
rect 666 19347 734 19403
rect 790 19347 858 19403
rect 914 19347 982 19403
rect 1038 19347 1106 19403
rect 1162 19347 1230 19403
rect 1286 19347 1354 19403
rect 1410 19347 1478 19403
rect 1534 19347 1602 19403
rect 1658 19347 1726 19403
rect 1782 19347 1850 19403
rect 1906 19347 2000 19403
rect 0 19279 2000 19347
rect 0 19223 114 19279
rect 170 19223 238 19279
rect 294 19223 362 19279
rect 418 19223 486 19279
rect 542 19223 610 19279
rect 666 19223 734 19279
rect 790 19223 858 19279
rect 914 19223 982 19279
rect 1038 19223 1106 19279
rect 1162 19223 1230 19279
rect 1286 19223 1354 19279
rect 1410 19223 1478 19279
rect 1534 19223 1602 19279
rect 1658 19223 1726 19279
rect 1782 19223 1850 19279
rect 1906 19223 2000 19279
rect 0 19155 2000 19223
rect 0 19099 114 19155
rect 170 19099 238 19155
rect 294 19099 362 19155
rect 418 19099 486 19155
rect 542 19099 610 19155
rect 666 19099 734 19155
rect 790 19099 858 19155
rect 914 19099 982 19155
rect 1038 19099 1106 19155
rect 1162 19099 1230 19155
rect 1286 19099 1354 19155
rect 1410 19099 1478 19155
rect 1534 19099 1602 19155
rect 1658 19099 1726 19155
rect 1782 19099 1850 19155
rect 1906 19099 2000 19155
rect 0 19031 2000 19099
rect 0 18975 114 19031
rect 170 18975 238 19031
rect 294 18975 362 19031
rect 418 18975 486 19031
rect 542 18975 610 19031
rect 666 18975 734 19031
rect 790 18975 858 19031
rect 914 18975 982 19031
rect 1038 18975 1106 19031
rect 1162 18975 1230 19031
rect 1286 18975 1354 19031
rect 1410 18975 1478 19031
rect 1534 18975 1602 19031
rect 1658 18975 1726 19031
rect 1782 18975 1850 19031
rect 1906 18975 2000 19031
rect 0 18907 2000 18975
rect 0 18851 114 18907
rect 170 18851 238 18907
rect 294 18851 362 18907
rect 418 18851 486 18907
rect 542 18851 610 18907
rect 666 18851 734 18907
rect 790 18851 858 18907
rect 914 18851 982 18907
rect 1038 18851 1106 18907
rect 1162 18851 1230 18907
rect 1286 18851 1354 18907
rect 1410 18851 1478 18907
rect 1534 18851 1602 18907
rect 1658 18851 1726 18907
rect 1782 18851 1850 18907
rect 1906 18851 2000 18907
rect 0 18783 2000 18851
rect 0 18727 114 18783
rect 170 18727 238 18783
rect 294 18727 362 18783
rect 418 18727 486 18783
rect 542 18727 610 18783
rect 666 18727 734 18783
rect 790 18727 858 18783
rect 914 18727 982 18783
rect 1038 18727 1106 18783
rect 1162 18727 1230 18783
rect 1286 18727 1354 18783
rect 1410 18727 1478 18783
rect 1534 18727 1602 18783
rect 1658 18727 1726 18783
rect 1782 18727 1850 18783
rect 1906 18727 2000 18783
rect 0 18659 2000 18727
rect 0 18603 114 18659
rect 170 18603 238 18659
rect 294 18603 362 18659
rect 418 18603 486 18659
rect 542 18603 610 18659
rect 666 18603 734 18659
rect 790 18603 858 18659
rect 914 18603 982 18659
rect 1038 18603 1106 18659
rect 1162 18603 1230 18659
rect 1286 18603 1354 18659
rect 1410 18603 1478 18659
rect 1534 18603 1602 18659
rect 1658 18603 1726 18659
rect 1782 18603 1850 18659
rect 1906 18603 2000 18659
rect 0 18535 2000 18603
rect 0 18479 114 18535
rect 170 18479 238 18535
rect 294 18479 362 18535
rect 418 18479 486 18535
rect 542 18479 610 18535
rect 666 18479 734 18535
rect 790 18479 858 18535
rect 914 18479 982 18535
rect 1038 18479 1106 18535
rect 1162 18479 1230 18535
rect 1286 18479 1354 18535
rect 1410 18479 1478 18535
rect 1534 18479 1602 18535
rect 1658 18479 1726 18535
rect 1782 18479 1850 18535
rect 1906 18479 2000 18535
rect 0 18411 2000 18479
rect 0 18355 114 18411
rect 170 18355 238 18411
rect 294 18355 362 18411
rect 418 18355 486 18411
rect 542 18355 610 18411
rect 666 18355 734 18411
rect 790 18355 858 18411
rect 914 18355 982 18411
rect 1038 18355 1106 18411
rect 1162 18355 1230 18411
rect 1286 18355 1354 18411
rect 1410 18355 1478 18411
rect 1534 18355 1602 18411
rect 1658 18355 1726 18411
rect 1782 18355 1850 18411
rect 1906 18355 2000 18411
rect 0 18287 2000 18355
rect 0 18231 114 18287
rect 170 18231 238 18287
rect 294 18231 362 18287
rect 418 18231 486 18287
rect 542 18231 610 18287
rect 666 18231 734 18287
rect 790 18231 858 18287
rect 914 18231 982 18287
rect 1038 18231 1106 18287
rect 1162 18231 1230 18287
rect 1286 18231 1354 18287
rect 1410 18231 1478 18287
rect 1534 18231 1602 18287
rect 1658 18231 1726 18287
rect 1782 18231 1850 18287
rect 1906 18231 2000 18287
rect 0 18163 2000 18231
rect 0 18107 114 18163
rect 170 18107 238 18163
rect 294 18107 362 18163
rect 418 18107 486 18163
rect 542 18107 610 18163
rect 666 18107 734 18163
rect 790 18107 858 18163
rect 914 18107 982 18163
rect 1038 18107 1106 18163
rect 1162 18107 1230 18163
rect 1286 18107 1354 18163
rect 1410 18107 1478 18163
rect 1534 18107 1602 18163
rect 1658 18107 1726 18163
rect 1782 18107 1850 18163
rect 1906 18107 2000 18163
rect 0 18039 2000 18107
rect 0 17983 114 18039
rect 170 17983 238 18039
rect 294 17983 362 18039
rect 418 17983 486 18039
rect 542 17983 610 18039
rect 666 17983 734 18039
rect 790 17983 858 18039
rect 914 17983 982 18039
rect 1038 17983 1106 18039
rect 1162 17983 1230 18039
rect 1286 17983 1354 18039
rect 1410 17983 1478 18039
rect 1534 17983 1602 18039
rect 1658 17983 1726 18039
rect 1782 17983 1850 18039
rect 1906 17983 2000 18039
rect 0 17915 2000 17983
rect 0 17859 114 17915
rect 170 17859 238 17915
rect 294 17859 362 17915
rect 418 17859 486 17915
rect 542 17859 610 17915
rect 666 17859 734 17915
rect 790 17859 858 17915
rect 914 17859 982 17915
rect 1038 17859 1106 17915
rect 1162 17859 1230 17915
rect 1286 17859 1354 17915
rect 1410 17859 1478 17915
rect 1534 17859 1602 17915
rect 1658 17859 1726 17915
rect 1782 17859 1850 17915
rect 1906 17859 2000 17915
rect 0 17791 2000 17859
rect 0 17735 114 17791
rect 170 17735 238 17791
rect 294 17735 362 17791
rect 418 17735 486 17791
rect 542 17735 610 17791
rect 666 17735 734 17791
rect 790 17735 858 17791
rect 914 17735 982 17791
rect 1038 17735 1106 17791
rect 1162 17735 1230 17791
rect 1286 17735 1354 17791
rect 1410 17735 1478 17791
rect 1534 17735 1602 17791
rect 1658 17735 1726 17791
rect 1782 17735 1850 17791
rect 1906 17735 2000 17791
rect 0 17667 2000 17735
rect 0 17611 114 17667
rect 170 17611 238 17667
rect 294 17611 362 17667
rect 418 17611 486 17667
rect 542 17611 610 17667
rect 666 17611 734 17667
rect 790 17611 858 17667
rect 914 17611 982 17667
rect 1038 17611 1106 17667
rect 1162 17611 1230 17667
rect 1286 17611 1354 17667
rect 1410 17611 1478 17667
rect 1534 17611 1602 17667
rect 1658 17611 1726 17667
rect 1782 17611 1850 17667
rect 1906 17611 2000 17667
rect 0 17543 2000 17611
rect 0 17487 114 17543
rect 170 17487 238 17543
rect 294 17487 362 17543
rect 418 17487 486 17543
rect 542 17487 610 17543
rect 666 17487 734 17543
rect 790 17487 858 17543
rect 914 17487 982 17543
rect 1038 17487 1106 17543
rect 1162 17487 1230 17543
rect 1286 17487 1354 17543
rect 1410 17487 1478 17543
rect 1534 17487 1602 17543
rect 1658 17487 1726 17543
rect 1782 17487 1850 17543
rect 1906 17487 2000 17543
rect 0 17419 2000 17487
rect 0 17363 114 17419
rect 170 17363 238 17419
rect 294 17363 362 17419
rect 418 17363 486 17419
rect 542 17363 610 17419
rect 666 17363 734 17419
rect 790 17363 858 17419
rect 914 17363 982 17419
rect 1038 17363 1106 17419
rect 1162 17363 1230 17419
rect 1286 17363 1354 17419
rect 1410 17363 1478 17419
rect 1534 17363 1602 17419
rect 1658 17363 1726 17419
rect 1782 17363 1850 17419
rect 1906 17363 2000 17419
rect 0 17200 2000 17363
rect 0 16852 2000 17000
rect 0 16796 114 16852
rect 170 16796 238 16852
rect 294 16796 362 16852
rect 418 16796 486 16852
rect 542 16796 610 16852
rect 666 16796 734 16852
rect 790 16796 858 16852
rect 914 16796 982 16852
rect 1038 16796 1106 16852
rect 1162 16796 1230 16852
rect 1286 16796 1354 16852
rect 1410 16796 1478 16852
rect 1534 16796 1602 16852
rect 1658 16796 1726 16852
rect 1782 16796 1850 16852
rect 1906 16796 2000 16852
rect 0 16728 2000 16796
rect 0 16672 114 16728
rect 170 16672 238 16728
rect 294 16672 362 16728
rect 418 16672 486 16728
rect 542 16672 610 16728
rect 666 16672 734 16728
rect 790 16672 858 16728
rect 914 16672 982 16728
rect 1038 16672 1106 16728
rect 1162 16672 1230 16728
rect 1286 16672 1354 16728
rect 1410 16672 1478 16728
rect 1534 16672 1602 16728
rect 1658 16672 1726 16728
rect 1782 16672 1850 16728
rect 1906 16672 2000 16728
rect 0 16604 2000 16672
rect 0 16548 114 16604
rect 170 16548 238 16604
rect 294 16548 362 16604
rect 418 16548 486 16604
rect 542 16548 610 16604
rect 666 16548 734 16604
rect 790 16548 858 16604
rect 914 16548 982 16604
rect 1038 16548 1106 16604
rect 1162 16548 1230 16604
rect 1286 16548 1354 16604
rect 1410 16548 1478 16604
rect 1534 16548 1602 16604
rect 1658 16548 1726 16604
rect 1782 16548 1850 16604
rect 1906 16548 2000 16604
rect 0 16480 2000 16548
rect 0 16424 114 16480
rect 170 16424 238 16480
rect 294 16424 362 16480
rect 418 16424 486 16480
rect 542 16424 610 16480
rect 666 16424 734 16480
rect 790 16424 858 16480
rect 914 16424 982 16480
rect 1038 16424 1106 16480
rect 1162 16424 1230 16480
rect 1286 16424 1354 16480
rect 1410 16424 1478 16480
rect 1534 16424 1602 16480
rect 1658 16424 1726 16480
rect 1782 16424 1850 16480
rect 1906 16424 2000 16480
rect 0 16356 2000 16424
rect 0 16300 114 16356
rect 170 16300 238 16356
rect 294 16300 362 16356
rect 418 16300 486 16356
rect 542 16300 610 16356
rect 666 16300 734 16356
rect 790 16300 858 16356
rect 914 16300 982 16356
rect 1038 16300 1106 16356
rect 1162 16300 1230 16356
rect 1286 16300 1354 16356
rect 1410 16300 1478 16356
rect 1534 16300 1602 16356
rect 1658 16300 1726 16356
rect 1782 16300 1850 16356
rect 1906 16300 2000 16356
rect 0 16232 2000 16300
rect 0 16176 114 16232
rect 170 16176 238 16232
rect 294 16176 362 16232
rect 418 16176 486 16232
rect 542 16176 610 16232
rect 666 16176 734 16232
rect 790 16176 858 16232
rect 914 16176 982 16232
rect 1038 16176 1106 16232
rect 1162 16176 1230 16232
rect 1286 16176 1354 16232
rect 1410 16176 1478 16232
rect 1534 16176 1602 16232
rect 1658 16176 1726 16232
rect 1782 16176 1850 16232
rect 1906 16176 2000 16232
rect 0 16108 2000 16176
rect 0 16052 114 16108
rect 170 16052 238 16108
rect 294 16052 362 16108
rect 418 16052 486 16108
rect 542 16052 610 16108
rect 666 16052 734 16108
rect 790 16052 858 16108
rect 914 16052 982 16108
rect 1038 16052 1106 16108
rect 1162 16052 1230 16108
rect 1286 16052 1354 16108
rect 1410 16052 1478 16108
rect 1534 16052 1602 16108
rect 1658 16052 1726 16108
rect 1782 16052 1850 16108
rect 1906 16052 2000 16108
rect 0 15984 2000 16052
rect 0 15928 114 15984
rect 170 15928 238 15984
rect 294 15928 362 15984
rect 418 15928 486 15984
rect 542 15928 610 15984
rect 666 15928 734 15984
rect 790 15928 858 15984
rect 914 15928 982 15984
rect 1038 15928 1106 15984
rect 1162 15928 1230 15984
rect 1286 15928 1354 15984
rect 1410 15928 1478 15984
rect 1534 15928 1602 15984
rect 1658 15928 1726 15984
rect 1782 15928 1850 15984
rect 1906 15928 2000 15984
rect 0 15860 2000 15928
rect 0 15804 114 15860
rect 170 15804 238 15860
rect 294 15804 362 15860
rect 418 15804 486 15860
rect 542 15804 610 15860
rect 666 15804 734 15860
rect 790 15804 858 15860
rect 914 15804 982 15860
rect 1038 15804 1106 15860
rect 1162 15804 1230 15860
rect 1286 15804 1354 15860
rect 1410 15804 1478 15860
rect 1534 15804 1602 15860
rect 1658 15804 1726 15860
rect 1782 15804 1850 15860
rect 1906 15804 2000 15860
rect 0 15736 2000 15804
rect 0 15680 114 15736
rect 170 15680 238 15736
rect 294 15680 362 15736
rect 418 15680 486 15736
rect 542 15680 610 15736
rect 666 15680 734 15736
rect 790 15680 858 15736
rect 914 15680 982 15736
rect 1038 15680 1106 15736
rect 1162 15680 1230 15736
rect 1286 15680 1354 15736
rect 1410 15680 1478 15736
rect 1534 15680 1602 15736
rect 1658 15680 1726 15736
rect 1782 15680 1850 15736
rect 1906 15680 2000 15736
rect 0 15612 2000 15680
rect 0 15556 114 15612
rect 170 15556 238 15612
rect 294 15556 362 15612
rect 418 15556 486 15612
rect 542 15556 610 15612
rect 666 15556 734 15612
rect 790 15556 858 15612
rect 914 15556 982 15612
rect 1038 15556 1106 15612
rect 1162 15556 1230 15612
rect 1286 15556 1354 15612
rect 1410 15556 1478 15612
rect 1534 15556 1602 15612
rect 1658 15556 1726 15612
rect 1782 15556 1850 15612
rect 1906 15556 2000 15612
rect 0 15488 2000 15556
rect 0 15432 114 15488
rect 170 15432 238 15488
rect 294 15432 362 15488
rect 418 15432 486 15488
rect 542 15432 610 15488
rect 666 15432 734 15488
rect 790 15432 858 15488
rect 914 15432 982 15488
rect 1038 15432 1106 15488
rect 1162 15432 1230 15488
rect 1286 15432 1354 15488
rect 1410 15432 1478 15488
rect 1534 15432 1602 15488
rect 1658 15432 1726 15488
rect 1782 15432 1850 15488
rect 1906 15432 2000 15488
rect 0 15364 2000 15432
rect 0 15308 114 15364
rect 170 15308 238 15364
rect 294 15308 362 15364
rect 418 15308 486 15364
rect 542 15308 610 15364
rect 666 15308 734 15364
rect 790 15308 858 15364
rect 914 15308 982 15364
rect 1038 15308 1106 15364
rect 1162 15308 1230 15364
rect 1286 15308 1354 15364
rect 1410 15308 1478 15364
rect 1534 15308 1602 15364
rect 1658 15308 1726 15364
rect 1782 15308 1850 15364
rect 1906 15308 2000 15364
rect 0 15240 2000 15308
rect 0 15184 114 15240
rect 170 15184 238 15240
rect 294 15184 362 15240
rect 418 15184 486 15240
rect 542 15184 610 15240
rect 666 15184 734 15240
rect 790 15184 858 15240
rect 914 15184 982 15240
rect 1038 15184 1106 15240
rect 1162 15184 1230 15240
rect 1286 15184 1354 15240
rect 1410 15184 1478 15240
rect 1534 15184 1602 15240
rect 1658 15184 1726 15240
rect 1782 15184 1850 15240
rect 1906 15184 2000 15240
rect 0 15116 2000 15184
rect 0 15060 114 15116
rect 170 15060 238 15116
rect 294 15060 362 15116
rect 418 15060 486 15116
rect 542 15060 610 15116
rect 666 15060 734 15116
rect 790 15060 858 15116
rect 914 15060 982 15116
rect 1038 15060 1106 15116
rect 1162 15060 1230 15116
rect 1286 15060 1354 15116
rect 1410 15060 1478 15116
rect 1534 15060 1602 15116
rect 1658 15060 1726 15116
rect 1782 15060 1850 15116
rect 1906 15060 2000 15116
rect 0 14992 2000 15060
rect 0 14936 114 14992
rect 170 14936 238 14992
rect 294 14936 362 14992
rect 418 14936 486 14992
rect 542 14936 610 14992
rect 666 14936 734 14992
rect 790 14936 858 14992
rect 914 14936 982 14992
rect 1038 14936 1106 14992
rect 1162 14936 1230 14992
rect 1286 14936 1354 14992
rect 1410 14936 1478 14992
rect 1534 14936 1602 14992
rect 1658 14936 1726 14992
rect 1782 14936 1850 14992
rect 1906 14936 2000 14992
rect 0 14868 2000 14936
rect 0 14812 114 14868
rect 170 14812 238 14868
rect 294 14812 362 14868
rect 418 14812 486 14868
rect 542 14812 610 14868
rect 666 14812 734 14868
rect 790 14812 858 14868
rect 914 14812 982 14868
rect 1038 14812 1106 14868
rect 1162 14812 1230 14868
rect 1286 14812 1354 14868
rect 1410 14812 1478 14868
rect 1534 14812 1602 14868
rect 1658 14812 1726 14868
rect 1782 14812 1850 14868
rect 1906 14812 2000 14868
rect 0 14744 2000 14812
rect 0 14688 114 14744
rect 170 14688 238 14744
rect 294 14688 362 14744
rect 418 14688 486 14744
rect 542 14688 610 14744
rect 666 14688 734 14744
rect 790 14688 858 14744
rect 914 14688 982 14744
rect 1038 14688 1106 14744
rect 1162 14688 1230 14744
rect 1286 14688 1354 14744
rect 1410 14688 1478 14744
rect 1534 14688 1602 14744
rect 1658 14688 1726 14744
rect 1782 14688 1850 14744
rect 1906 14688 2000 14744
rect 0 14620 2000 14688
rect 0 14564 114 14620
rect 170 14564 238 14620
rect 294 14564 362 14620
rect 418 14564 486 14620
rect 542 14564 610 14620
rect 666 14564 734 14620
rect 790 14564 858 14620
rect 914 14564 982 14620
rect 1038 14564 1106 14620
rect 1162 14564 1230 14620
rect 1286 14564 1354 14620
rect 1410 14564 1478 14620
rect 1534 14564 1602 14620
rect 1658 14564 1726 14620
rect 1782 14564 1850 14620
rect 1906 14564 2000 14620
rect 0 14496 2000 14564
rect 0 14440 114 14496
rect 170 14440 238 14496
rect 294 14440 362 14496
rect 418 14440 486 14496
rect 542 14440 610 14496
rect 666 14440 734 14496
rect 790 14440 858 14496
rect 914 14440 982 14496
rect 1038 14440 1106 14496
rect 1162 14440 1230 14496
rect 1286 14440 1354 14496
rect 1410 14440 1478 14496
rect 1534 14440 1602 14496
rect 1658 14440 1726 14496
rect 1782 14440 1850 14496
rect 1906 14440 2000 14496
rect 0 14372 2000 14440
rect 0 14316 114 14372
rect 170 14316 238 14372
rect 294 14316 362 14372
rect 418 14316 486 14372
rect 542 14316 610 14372
rect 666 14316 734 14372
rect 790 14316 858 14372
rect 914 14316 982 14372
rect 1038 14316 1106 14372
rect 1162 14316 1230 14372
rect 1286 14316 1354 14372
rect 1410 14316 1478 14372
rect 1534 14316 1602 14372
rect 1658 14316 1726 14372
rect 1782 14316 1850 14372
rect 1906 14316 2000 14372
rect 0 14248 2000 14316
rect 0 14192 114 14248
rect 170 14192 238 14248
rect 294 14192 362 14248
rect 418 14192 486 14248
rect 542 14192 610 14248
rect 666 14192 734 14248
rect 790 14192 858 14248
rect 914 14192 982 14248
rect 1038 14192 1106 14248
rect 1162 14192 1230 14248
rect 1286 14192 1354 14248
rect 1410 14192 1478 14248
rect 1534 14192 1602 14248
rect 1658 14192 1726 14248
rect 1782 14192 1850 14248
rect 1906 14192 2000 14248
rect 0 14000 2000 14192
use GF_NI_FILL10_1short  GF_NI_FILL10_1_0
timestamp 1765934810
transform 1 0 0 0 1 0
box -32 13097 2032 69968
<< labels >>
rlabel metal4 s 1018 18921 1018 18921 4 DVSS
port 1 nsew
rlabel metal4 s 1018 15750 1018 15750 4 DVSS
port 1 nsew
rlabel metal4 s 1018 21907 1018 21907 4 DVSS
port 1 nsew
rlabel metal4 s 1018 26100 1018 26100 4 DVSS
port 1 nsew
rlabel metal4 s 1018 40342 1018 40342 4 DVSS
port 1 nsew
rlabel metal4 s 1018 47595 1018 47595 4 DVSS
port 1 nsew
rlabel metal4 s 1018 57858 1018 57858 4 DVSS
port 1 nsew
rlabel metal4 s 1018 61058 1018 61058 4 DVSS
port 1 nsew
rlabel metal4 s 1018 66023 1018 66023 4 DVSS
port 1 nsew
rlabel metal4 s 1018 69049 1018 69049 4 DVSS
port 1 nsew
rlabel metal3 s 1018 69049 1018 69049 4 DVSS
port 1 nsew
rlabel metal3 s 1018 40342 1018 40342 4 DVSS
port 1 nsew
rlabel metal3 s 1018 26100 1018 26100 4 DVSS
port 1 nsew
rlabel metal3 s 1018 21907 1018 21907 4 DVSS
port 1 nsew
rlabel metal3 s 1018 18921 1018 18921 4 DVSS
port 1 nsew
rlabel metal3 s 1018 15750 1018 15750 4 DVSS
port 1 nsew
rlabel metal3 s 1018 61058 1018 61058 4 DVSS
port 1 nsew
rlabel metal3 s 1018 57858 1018 57858 4 DVSS
port 1 nsew
rlabel metal3 s 1018 47595 1018 47595 4 DVSS
port 1 nsew
rlabel metal3 s 1018 66023 1018 66023 4 DVSS
port 1 nsew
rlabel metal4 s 1018 31609 1018 31609 4 DVDD
port 2 nsew
rlabel metal4 s 1018 28394 1018 28394 4 DVDD
port 2 nsew
rlabel metal4 s 1018 24284 1018 24284 4 DVDD
port 2 nsew
rlabel metal4 s 1018 59623 1018 59623 4 DVDD
port 2 nsew
rlabel metal4 s 1018 56423 1018 56423 4 DVDD
port 2 nsew
rlabel metal4 s 1018 54658 1018 54658 4 DVDD
port 2 nsew
rlabel metal4 s 1018 53223 1018 53223 4 DVDD
port 2 nsew
rlabel metal4 s 1018 44368 1018 44368 4 DVDD
port 2 nsew
rlabel metal4 s 1018 41977 1018 41977 4 DVDD
port 2 nsew
rlabel metal4 s 1018 37959 1018 37959 4 DVDD
port 2 nsew
rlabel metal4 s 1018 34723 1018 34723 4 DVDD
port 2 nsew
rlabel metal4 s 1018 67458 1018 67458 4 DVDD
port 2 nsew
rlabel metal3 s 1018 41977 1018 41977 4 DVDD
port 2 nsew
rlabel metal3 s 1018 37959 1018 37959 4 DVDD
port 2 nsew
rlabel metal3 s 1018 34723 1018 34723 4 DVDD
port 2 nsew
rlabel metal3 s 1018 31609 1018 31609 4 DVDD
port 2 nsew
rlabel metal3 s 1018 28394 1018 28394 4 DVDD
port 2 nsew
rlabel metal3 s 1018 24284 1018 24284 4 DVDD
port 2 nsew
rlabel metal3 s 1018 59623 1018 59623 4 DVDD
port 2 nsew
rlabel metal3 s 1018 56423 1018 56423 4 DVDD
port 2 nsew
rlabel metal3 s 1018 54658 1018 54658 4 DVDD
port 2 nsew
rlabel metal3 s 1018 53223 1018 53223 4 DVDD
port 2 nsew
rlabel metal3 s 1018 44368 1018 44368 4 DVDD
port 2 nsew
rlabel metal3 s 1018 67458 1018 67458 4 DVDD
port 2 nsew
rlabel metal4 s 1018 51458 1018 51458 4 VDD
port 3 nsew
rlabel metal4 s 1018 62823 1018 62823 4 VDD
port 3 nsew
rlabel metal3 s 1018 51458 1018 51458 4 VDD
port 3 nsew
rlabel metal3 s 1018 62823 1018 62823 4 VDD
port 3 nsew
rlabel metal4 s 1018 64258 1018 64258 4 VSS
port 4 nsew
rlabel metal4 s 1018 50023 1018 50023 4 VSS
port 4 nsew
rlabel metal3 s 1018 50023 1018 50023 4 VSS
port 4 nsew
rlabel metal3 s 1018 64258 1018 64258 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2000 70000
<< end >>
