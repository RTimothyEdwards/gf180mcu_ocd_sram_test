magic
tech gf180mcuD
magscale 1 10
timestamp 1765233513
<< metal1 >>
rect 468012 150003 468673 150123
rect 468012 149219 468673 149339
<< via1 >>
rect 468981 149611 469040 149771
rect 469364 149608 469423 149768
rect 469485 149608 469544 149768
rect 470057 149632 470116 149792
rect 470885 149611 470944 149771
rect 471268 149608 471327 149768
rect 471389 149608 471448 149768
rect 471961 149632 472020 149792
rect 472789 149611 472848 149771
rect 473172 149608 473231 149768
rect 473293 149608 473352 149768
rect 473865 149632 473924 149792
rect 474693 149611 474752 149771
rect 475076 149608 475135 149768
rect 475197 149608 475256 149768
rect 475769 149632 475828 149792
rect 476597 149611 476656 149771
rect 476980 149608 477039 149768
rect 477101 149608 477160 149768
rect 477673 149632 477732 149792
rect 478501 149611 478560 149771
rect 478884 149608 478943 149768
rect 479005 149608 479064 149768
rect 479577 149632 479636 149792
rect 480405 149611 480464 149771
rect 480788 149608 480847 149768
rect 480909 149608 480968 149768
rect 481481 149632 481540 149792
rect 482309 149611 482368 149771
rect 482692 149608 482751 149768
rect 482813 149608 482872 149768
rect 483385 149632 483444 149792
<< metal2 >>
rect 469394 150646 469470 151238
rect 469394 150581 470119 150646
rect 468978 149771 469043 149790
rect 468978 149611 468981 149771
rect 469040 149611 469043 149771
rect 468978 148869 469043 149611
rect 469361 149768 469426 150336
rect 470054 149792 470119 150581
rect 471394 150598 471470 151238
rect 473394 150628 473470 151238
rect 471394 150548 472023 150598
rect 473394 150563 473927 150628
rect 471395 150533 472023 150548
rect 469361 149608 469364 149768
rect 469423 149608 469426 149768
rect 469361 149593 469426 149608
rect 469482 149768 469547 149787
rect 469482 149608 469485 149768
rect 469544 149608 469547 149768
rect 470054 149632 470057 149792
rect 470116 149632 470119 149792
rect 470054 149617 470119 149632
rect 470882 149771 470947 149790
rect 469482 148869 469547 149608
rect 470882 149611 470885 149771
rect 470944 149611 470947 149771
rect 470882 148869 470947 149611
rect 471265 149768 471330 150336
rect 471958 149792 472023 150533
rect 471265 149608 471268 149768
rect 471327 149608 471330 149768
rect 471265 149593 471330 149608
rect 471386 149768 471451 149787
rect 471386 149608 471389 149768
rect 471448 149608 471451 149768
rect 471958 149632 471961 149792
rect 472020 149632 472023 149792
rect 471958 149617 472023 149632
rect 472786 149771 472851 149790
rect 471386 148869 471451 149608
rect 472786 149611 472789 149771
rect 472848 149611 472851 149771
rect 472786 148869 472851 149611
rect 473169 149768 473234 150336
rect 473862 149792 473927 150563
rect 475394 150615 475470 151238
rect 475394 150550 475831 150615
rect 473169 149608 473172 149768
rect 473231 149608 473234 149768
rect 473169 149593 473234 149608
rect 473290 149768 473355 149787
rect 473290 149608 473293 149768
rect 473352 149608 473355 149768
rect 473862 149632 473865 149792
rect 473924 149632 473927 149792
rect 473862 149617 473927 149632
rect 474690 149771 474755 149790
rect 473290 148869 473355 149608
rect 474690 149611 474693 149771
rect 474752 149611 474755 149771
rect 474690 148869 474755 149611
rect 475073 149768 475138 150336
rect 475766 149792 475831 150550
rect 477394 150579 477470 151238
rect 479394 150590 479470 151238
rect 477394 150514 477735 150579
rect 479394 150525 479639 150590
rect 481394 150589 481470 151238
rect 483394 150645 483470 151238
rect 475073 149608 475076 149768
rect 475135 149608 475138 149768
rect 475073 149593 475138 149608
rect 475194 149768 475259 149787
rect 475194 149608 475197 149768
rect 475256 149608 475259 149768
rect 475766 149632 475769 149792
rect 475828 149632 475831 149792
rect 475766 149617 475831 149632
rect 476594 149771 476659 149790
rect 475194 148869 475259 149608
rect 476594 149611 476597 149771
rect 476656 149611 476659 149771
rect 476594 148869 476659 149611
rect 476977 149768 477042 150336
rect 477670 149792 477735 150514
rect 476977 149608 476980 149768
rect 477039 149608 477042 149768
rect 476977 149593 477042 149608
rect 477098 149768 477163 149787
rect 477098 149608 477101 149768
rect 477160 149608 477163 149768
rect 477670 149632 477673 149792
rect 477732 149632 477735 149792
rect 477670 149617 477735 149632
rect 478498 149771 478563 149790
rect 477098 148869 477163 149608
rect 478498 149611 478501 149771
rect 478560 149611 478563 149771
rect 478498 148869 478563 149611
rect 478881 149768 478946 150336
rect 479574 149792 479639 150525
rect 481393 150524 481543 150589
rect 478881 149608 478884 149768
rect 478943 149608 478946 149768
rect 478881 149593 478946 149608
rect 479002 149768 479067 149787
rect 479002 149608 479005 149768
rect 479064 149608 479067 149768
rect 479574 149632 479577 149792
rect 479636 149632 479639 149792
rect 479574 149617 479639 149632
rect 480402 149771 480467 149790
rect 479002 148869 479067 149608
rect 480402 149611 480405 149771
rect 480464 149611 480467 149771
rect 480402 148869 480467 149611
rect 480785 149768 480850 150336
rect 481478 149792 481543 150524
rect 483382 150548 483470 150645
rect 480785 149608 480788 149768
rect 480847 149608 480850 149768
rect 480785 149593 480850 149608
rect 480906 149768 480971 149787
rect 480906 149608 480909 149768
rect 480968 149608 480971 149768
rect 481478 149632 481481 149792
rect 481540 149632 481543 149792
rect 481478 149617 481543 149632
rect 482306 149771 482371 149790
rect 480906 148869 480971 149608
rect 482306 149611 482309 149771
rect 482368 149611 482371 149771
rect 482306 148869 482371 149611
rect 482689 149768 482754 150336
rect 483382 149792 483447 150548
rect 482689 149608 482692 149768
rect 482751 149608 482754 149768
rect 482689 149593 482754 149608
rect 482810 149768 482875 149787
rect 482810 149608 482813 149768
rect 482872 149608 482875 149768
rect 483382 149632 483385 149792
rect 483444 149632 483447 149792
rect 483382 149617 483447 149632
rect 482810 148869 482875 149608
<< metal3 >>
rect 467911 150270 483680 150346
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_2 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 468012 0 1 149279
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_3
timestamp 1751532246
transform 1 0 483916 0 1 149279
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_8 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914320
transform 1 0 470588 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_9
timestamp 1751914320
transform 1 0 468684 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_10
timestamp 1751914320
transform 1 0 476300 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_11
timestamp 1751914320
transform 1 0 474396 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_12
timestamp 1751914320
transform 1 0 472492 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_13
timestamp 1751914320
transform 1 0 482012 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_14
timestamp 1751914320
transform 1 0 480108 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__mux2_4  gf180mcu_as_sc_mcu7t3v3__mux2_4_15
timestamp 1751914320
transform 1 0 478204 0 1 149279
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_9 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1759751540
transform 1 0 468460 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_10
timestamp 1759751540
transform 1 0 470364 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_11
timestamp 1759751540
transform 1 0 476076 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_12
timestamp 1759751540
transform 1 0 474172 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_13
timestamp 1759751540
transform 1 0 472268 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_14
timestamp 1759751540
transform 1 0 483692 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_15
timestamp 1759751540
transform 1 0 481788 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_16
timestamp 1759751540
transform 1 0 479884 0 1 149279
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_17
timestamp 1759751540
transform 1 0 477980 0 1 149279
box -86 -86 310 870
use ocd_via2_3x  ocd_via2_3x_229
timestamp 1765059587
transform 1 0 381396 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_230
timestamp 1765059587
transform 1 0 379492 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_231
timestamp 1765059587
transform 1 0 387108 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_232
timestamp 1765059587
transform 1 0 385204 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_233
timestamp 1765059587
transform 1 0 383300 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_234
timestamp 1765059587
transform 1 0 392820 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_235
timestamp 1765059587
transform 1 0 390916 0 1 3830
box 89752 146428 90065 146528
use ocd_via2_3x  ocd_via2_3x_236
timestamp 1765059587
transform 1 0 389012 0 1 3830
box 89752 146428 90065 146528
<< labels >>
flabel metal1 468012 150003 468673 150123 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal1 468012 149219 468673 149339 0 FreeSans 480 0 0 0 vss
port 1 nsew
flabel metal3 467911 150270 468070 150346 0 FreeSans 480 0 0 0 S
port 2 nsew
flabel metal2 469482 148869 469547 148932 0 FreeSans 480 0 0 0 A[7]
port 3 nsew
flabel metal2 471386 148869 471451 148932 0 FreeSans 480 0 0 0 A[6]
port 4 nsew
flabel metal2 473290 148869 473355 148932 0 FreeSans 480 0 0 0 A[5]
port 5 nsew
flabel metal2 475194 148869 475259 148932 0 FreeSans 480 0 0 0 A[4]
port 6 nsew
flabel metal2 477098 148869 477163 148932 0 FreeSans 480 0 0 0 A[3]
port 7 nsew
flabel metal2 479002 148869 479067 148932 0 FreeSans 480 0 0 0 A[2]
port 8 nsew
flabel metal2 480906 148869 480971 148932 0 FreeSans 480 0 0 0 A[1]
port 9 nsew
flabel metal2 482810 148869 482875 148932 0 FreeSans 480 0 0 0 A[0]
port 10 nsew
flabel metal2 468978 148869 469043 148932 0 FreeSans 480 0 0 0 B[7]
port 11 nsew
flabel metal2 470882 148869 470947 148932 0 FreeSans 480 0 0 0 B[6]
port 12 nsew
flabel metal2 472786 148869 472851 148932 0 FreeSans 480 0 0 0 B[5]
port 13 nsew
flabel metal2 474690 148869 474755 148932 0 FreeSans 480 0 0 0 B[4]
port 14 nsew
flabel metal2 476594 148869 476659 148932 0 FreeSans 480 0 0 0 B[3]
port 15 nsew
flabel metal2 478498 148869 478563 148932 0 FreeSans 480 0 0 0 B[2]
port 16 nsew
flabel metal2 480402 148869 480467 148932 0 FreeSans 480 0 0 0 B[1]
port 17 nsew
flabel metal2 482306 148869 482371 148932 0 FreeSans 480 0 0 0 B[0]
port 18 nsew
flabel metal2 469394 151166 469470 151238 0 FreeSans 480 0 0 0 Y[7]
port 19 nsew
flabel metal2 471394 151166 471470 151238 0 FreeSans 480 0 0 0 Y[6]
port 20 nsew
flabel metal2 473394 151166 473470 151238 0 FreeSans 480 0 0 0 Y[5]
port 21 nsew
flabel metal2 475394 151166 475470 151238 0 FreeSans 480 0 0 0 Y[4]
port 22 nsew
flabel metal2 477394 151166 477470 151238 0 FreeSans 480 0 0 0 Y[3]
port 23 nsew
flabel metal2 479394 151166 479470 151238 0 FreeSans 480 0 0 0 Y[2]
port 24 nsew
flabel metal2 481394 151166 481470 151238 0 FreeSans 480 0 0 0 Y[1]
port 25 nsew
flabel metal2 483394 151166 483470 151238 0 FreeSans 480 0 0 0 Y[0]
port 26 nsew
<< end >>
