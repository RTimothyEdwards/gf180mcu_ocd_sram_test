magic
tech gf180mcuD
magscale 1 10
timestamp 1765054368
<< metal1 >>
rect 0 133 14889 185
rect 15055 133 15452 185
rect 0 35 15345 87
rect 15511 35 15527 87
<< via1 >>
rect 14889 133 15055 185
rect 15345 35 15511 87
<< metal2 >>
rect 182 -48 258 232
rect 703 -48 779 232
rect 932 -48 1008 232
rect 1074 -48 1150 232
rect 1216 -48 1292 232
rect 1576 -48 1652 232
rect 1787 -48 1863 232
rect 13244 -48 13320 232
rect 13390 -48 13466 232
rect 13536 -48 13612 232
rect 13682 -48 13758 232
rect 15068 187 15144 232
rect 14877 185 15144 187
rect 14877 133 14889 185
rect 15055 133 15144 185
rect 14877 131 15144 133
rect 15068 0 15144 131
rect 15256 89 15332 232
rect 15256 87 15523 89
rect 15256 35 15345 87
rect 15511 35 15523 87
rect 15256 33 15523 35
rect 15256 0 15332 33
<< end >>
