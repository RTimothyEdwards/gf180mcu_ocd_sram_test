* NGSPICE file created from gf180mcu_ocd_sram_test.ext - technology: gf180mcuD

.subckt pmos_5p04310591302061_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1836p pd=6.26u as=1.1836p ps=6.26u w=2.69u l=0.28u
.ends

.subckt pmos_1p2$$47820844_3v512x8m81 a_n14_n34# pmos_5p04310591302061_3v512x8m81_0/S
+ w_n133_n65# pmos_5p04310591302061_3v512x8m81_0/D
Xpmos_5p04310591302061_3v512x8m81_0 pmos_5p04310591302061_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302061_3v512x8m81_0/S pmos_5p04310591302061_3v512x8m81
.ends

.subckt pmos_5p04310591302060_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1638p pd=6.17u as=1.1638p ps=6.17u w=2.645u l=0.28u
.ends

.subckt pmos_1p2$$47821868_3v512x8m81 pmos_5p04310591302060_3v512x8m81_0/S w_n133_n66#
+ a_n14_n34# pmos_5p04310591302060_3v512x8m81_0/D
Xpmos_5p04310591302060_3v512x8m81_0 pmos_5p04310591302060_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302060_3v512x8m81_0/S pmos_5p04310591302060_3v512x8m81
.ends

.subckt nmos_5p04310591302010_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$46551084_3v512x8m81 nmos_5p04310591302010_3v512x8m81_0/S nmos_5p04310591302010_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302010_3v512x8m81_0 nmos_5p04310591302010_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v512x8m81_0/S VSUBS nmos_5p04310591302010_3v512x8m81
.ends

.subckt ypredec1_xa_3v512x8m81 m1_n40_n2861# pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_145_n4683# m3_0_n4986# m1_n40_n3567# m1_n40_n3285# a_0_56# pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_465_n4683# M2_M1$$47515692_3v512x8m81_0/VSUBS m1_n40_n3426# m1_n40_n3144# m1_n40_n3003#
+ a_305_n4683# pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
Xpmos_1p2$$47820844_3v512x8m81_0 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D pmos_1p2$$47820844_3v512x8m81
Xpmos_1p2$$47820844_3v512x8m81_1 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S pmos_1p2$$47820844_3v512x8m81
Xpmos_1p2$$47820844_3v512x8m81_2 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D pmos_1p2$$47820844_3v512x8m81
Xpmos_1p2$$47821868_3v512x8m81_0 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66# a_145_n4683# pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81
Xnmos_1p2$$46551084_3v512x8m81_0 pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M2_M1$$47515692_3v512x8m81_0/VSUBS pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ M2_M1$$47515692_3v512x8m81_0/VSUBS nmos_1p2$$46551084_3v512x8m81
Xnmos_1p2$$46551084_3v512x8m81_1 M2_M1$$47515692_3v512x8m81_0/VSUBS pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D M2_M1$$47515692_3v512x8m81_0/VSUBS
+ nmos_1p2$$46551084_3v512x8m81
Xpmos_1p2$$47821868_3v512x8m81_2 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66# a_305_n4683# pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ pmos_1p2$$47821868_3v512x8m81
Xnmos_1p2$$46551084_3v512x8m81_2 M2_M1$$47515692_3v512x8m81_0/VSUBS pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D M2_M1$$47515692_3v512x8m81_0/VSUBS
+ nmos_1p2$$46551084_3v512x8m81
Xpmos_1p2$$47821868_3v512x8m81_3 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66# a_465_n4683# pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D
+ pmos_1p2$$47821868_3v512x8m81
X0 a_361_n4624# a_305_n4683# a_201_n4624# M2_M1$$47515692_3v512x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=0.8268p ps=3.7u w=3.18u l=0.28u
X1 a_201_n4624# a_145_n4683# M2_M1$$47515692_3v512x8m81_0/VSUBS M2_M1$$47515692_3v512x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=1.4469p ps=7.27u w=3.18u l=0.28u
X2 pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/D a_465_n4683# a_361_n4624# M2_M1$$47515692_3v512x8m81_0/VSUBS nfet_03v3 ad=1.5423p pd=7.33u as=0.8268p ps=3.7u w=3.18u l=0.28u
.ends

.subckt ypredec1_xax8_3v512x8m81 ypredec1_xa_3v512x8m81_0/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xa_3v512x8m81_5/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_997_2070# ypredec1_xa_3v512x8m81_1/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xa_3v512x8m81_6/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xa_3v512x8m81_5/a_0_56# ypredec1_xa_3v512x8m81_2/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_683_1364# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_4427_1646# ypredec1_xa_3v512x8m81_3/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_4270_1505# a_526_1788# ypredec1_xa_3v512x8m81_3/a_0_56# ypredec1_xa_3v512x8m81_4/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_840_1930# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ VSUBS ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
Xypredec1_xa_3v512x8m81_0 a_997_2070# ypredec1_xa_3v512x8m81_0/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_0/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_4427_1646# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_840_1930# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_1 a_997_2070# ypredec1_xa_3v512x8m81_1/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_5/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_4427_1646# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_4270_1505# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_2 a_997_2070# ypredec1_xa_3v512x8m81_2/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_526_1788# VSUBS a_683_1364# a_4427_1646# VSUBS ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_997_2070# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_4270_1505# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_3 a_997_2070# ypredec1_xa_3v512x8m81_3/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_3/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_997_2070# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_840_1930# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_4 a_997_2070# ypredec1_xa_3v512x8m81_4/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_4/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_4427_1646# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_840_1930# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_5 a_997_2070# ypredec1_xa_3v512x8m81_5/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_5/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_4427_1646# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_4270_1505# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_6 a_997_2070# ypredec1_xa_3v512x8m81_6/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_6/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_997_2070# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_4270_1505# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
Xypredec1_xa_3v512x8m81_7 a_997_2070# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v512x8m81_7/a_0_56# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/w_n133_n65#
+ a_997_2070# VSUBS a_4270_1505# a_526_1788# a_840_1930# a_840_1930# ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/w_n133_n66#
+ ypredec1_xa_3v512x8m81_7/pmos_1p2$$47821868_3v512x8m81_3/pmos_5p04310591302060_3v512x8m81_0/S
+ ypredec1_xa_3v512x8m81
.ends

.subckt pmos_5p04310591302055_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.1052p pd=19.54u as=4.1052p ps=19.54u w=9.33u l=0.28u
.ends

.subckt nmos_5p04310591302054_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.8634p pd=9.35u as=1.8634p ps=9.35u w=4.235u l=0.28u
.ends

.subckt ypredec1_ys_3v512x8m81 a_161_1551# nmos_5p04310591302054_3v512x8m81_1/D pmos_5p04310591302055_3v512x8m81_1/S
+ nmos_5p04310591302054_3v512x8m81_3/D nmos_5p04310591302054_3v512x8m81_2/S pmos_5p04310591302055_3v512x8m81_3/S
+ pmos_5p04310591302055_3v512x8m81_3/D VSUBS
Xpmos_5p04310591302055_3v512x8m81_2 pmos_5p04310591302055_3v512x8m81_3/S pmos_5p04310591302055_3v512x8m81_0/D
+ pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81
Xpmos_5p04310591302055_3v512x8m81_3 pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_0/D
+ pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_3/S pmos_5p04310591302055_3v512x8m81
Xnmos_5p04310591302054_3v512x8m81_0 pmos_5p04310591302055_3v512x8m81_3/S pmos_5p04310591302055_3v512x8m81_0/D
+ nmos_5p04310591302054_3v512x8m81_1/D VSUBS nmos_5p04310591302054_3v512x8m81
Xnmos_5p04310591302054_3v512x8m81_1 nmos_5p04310591302054_3v512x8m81_1/D pmos_5p04310591302055_3v512x8m81_0/D
+ pmos_5p04310591302055_3v512x8m81_1/S VSUBS nmos_5p04310591302054_3v512x8m81
Xnmos_5p04310591302054_3v512x8m81_2 pmos_5p04310591302055_3v512x8m81_0/D a_161_1551#
+ nmos_5p04310591302054_3v512x8m81_2/S VSUBS nmos_5p04310591302054_3v512x8m81
Xnmos_5p04310591302054_3v512x8m81_3 nmos_5p04310591302054_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_0/D
+ pmos_5p04310591302055_3v512x8m81_3/S VSUBS nmos_5p04310591302054_3v512x8m81
Xpmos_5p04310591302055_3v512x8m81_0 pmos_5p04310591302055_3v512x8m81_0/D a_161_1551#
+ pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81
Xpmos_5p04310591302055_3v512x8m81_1 pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_0/D
+ pmos_5p04310591302055_3v512x8m81_3/D pmos_5p04310591302055_3v512x8m81_1/S pmos_5p04310591302055_3v512x8m81
.ends

.subckt pmos_5p04310591302062_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$47109164_3v512x8m81 pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ pmos_5p04310591302062_3v512x8m81_0/D a_118_159# pmos_5p04310591302062_3v512x8m81_0/S
+ a_n42_159#
Xpmos_5p04310591302062_3v512x8m81_0 pmos_5p04310591302062_3v512x8m81_0/D a_n42_159#
+ a_118_159# pmos_5p04310591302062_3v512x8m81_0/w_n202_n86# pmos_5p04310591302062_3v512x8m81_0/S
+ pmos_5p04310591302062_3v512x8m81
.ends

.subckt nmos_5p04310591302057_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.9306p pd=5.11u as=0.9306p ps=5.11u w=2.115u l=0.28u
.ends

.subckt nmos_1p2$$47514668_3v512x8m81 nmos_5p04310591302057_3v512x8m81_0/S nmos_5p04310591302057_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v512x8m81_0 nmos_5p04310591302057_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v512x8m81_0/S VSUBS nmos_5p04310591302057_3v512x8m81
.ends

.subckt pmos_5p0431059130204_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt pmos_1p2$$46887980_3v512x8m81 w_n133_n66# pmos_5p0431059130204_3v512x8m81_0/S
+ a_n14_n34# pmos_5p0431059130204_3v512x8m81_0/D
Xpmos_5p0431059130204_3v512x8m81_0 pmos_5p0431059130204_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130204_3v512x8m81_0/S pmos_5p0431059130204_3v512x8m81
.ends

.subckt nmos_5p04310591302059_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.28u
.ends

.subckt nmos_1p2$$47329324_3v512x8m81 nmos_5p04310591302059_3v512x8m81_0/D a_118_n34#
+ a_n41_n34# nmos_5p04310591302059_3v512x8m81_0/S VSUBS
Xnmos_5p04310591302059_3v512x8m81_0 nmos_5p04310591302059_3v512x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302059_3v512x8m81_0/S VSUBS nmos_5p04310591302059_3v512x8m81
.ends

.subckt pmos_5p04310591302041_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt pmos_1p2_161_3v512x8m81 pmos_5p04310591302041_3v512x8m81_0/D a_n14_89# pmos_5p04310591302041_3v512x8m81_0/S
+ w_n133_n65#
Xpmos_5p04310591302041_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81
.ends

.subckt nmos_1p2_157_3v512x8m81 nmos_5p04310591302010_3v512x8m81_0/S nmos_5p04310591302010_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302010_3v512x8m81_0 nmos_5p04310591302010_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v512x8m81_0/S VSUBS nmos_5p04310591302010_3v512x8m81
.ends

.subckt pmos_5p04310591302058_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.9306p pd=5.11u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$47331372_3v512x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302058_3v512x8m81_0/D
+ pmos_5p04310591302058_3v512x8m81_0/S a_118_n34#
Xpmos_5p04310591302058_3v512x8m81_0 pmos_5p04310591302058_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302058_3v512x8m81_0/S pmos_5p04310591302058_3v512x8m81
.ends

.subckt pmos_5p04310591302014_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2_160_3v512x8m81 w_n133_n66# pmos_5p04310591302014_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v512x8m81_0/D
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt alatch_3v512x8m81 enb en ab a vss a_886_665# vdd
Xnmos_1p2$$47329324_3v512x8m81_0 ab pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S vss vss nmos_1p2$$47329324_3v512x8m81
Xpmos_1p2_161_3v512x8m81_0 pmos_1p2_161_3v512x8m81_1/pmos_5p04310591302041_3v512x8m81_0/S
+ a_886_665# pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S vdd pmos_1p2_161_3v512x8m81
Xpmos_1p2_161_3v512x8m81_1 vdd ab pmos_1p2_161_3v512x8m81_1/pmos_5p04310591302041_3v512x8m81_0/S
+ vdd pmos_1p2_161_3v512x8m81
Xnmos_1p2_157_3v512x8m81_0 pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ a a_886_665# vss nmos_1p2_157_3v512x8m81
Xpmos_1p2$$47331372_3v512x8m81_0 pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ vdd ab vdd pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S pmos_1p2$$47331372_3v512x8m81
Xpmos_1p2_160_3v512x8m81_0 vdd pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ enb a pmos_1p2_160_3v512x8m81
X0 pmos_1p2_161_3v512x8m81_1/pmos_5p04310591302041_3v512x8m81_0/S enb pmos_1p2_161_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss ab pmos_1p2_161_3v512x8m81_1/pmos_5p04310591302041_3v512x8m81_0/S vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt ypredec1_bot_3v512x8m81 m1_n9_2295# m1_n9_2436# m1_n9_2154# m1_n9_2013# alatch_3v512x8m81_0/a
+ m1_n9_1871# pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ m1_n9_1730# pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ alatch_3v512x8m81_0/vss alatch_3v512x8m81_0/enb pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ m2_800_896# alatch_3v512x8m81_0/vdd
Xnmos_1p2$$47514668_3v512x8m81_0 alatch_3v512x8m81_0/vss pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D alatch_3v512x8m81_0/vss
+ nmos_1p2$$47514668_3v512x8m81
Xnmos_1p2$$47514668_3v512x8m81_1 alatch_3v512x8m81_0/vss pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ alatch_3v512x8m81_0/ab alatch_3v512x8m81_0/vss nmos_1p2$$47514668_3v512x8m81
Xpmos_1p2$$46887980_3v512x8m81_0 pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D pmos_1p2$$46887980_3v512x8m81
Xpmos_1p2$$46887980_3v512x8m81_1 pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S alatch_3v512x8m81_0/ab
+ pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D pmos_1p2$$46887980_3v512x8m81
Xalatch_3v512x8m81_0 alatch_3v512x8m81_0/enb alatch_3v512x8m81_0/en alatch_3v512x8m81_0/ab
+ alatch_3v512x8m81_0/a alatch_3v512x8m81_0/vss m2_800_896# alatch_3v512x8m81_0/vdd
+ alatch_3v512x8m81
.ends

.subckt nmos_5p04310591302056_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3916p pd=2.66u as=0.3916p ps=2.66u w=0.89u l=0.28u
.ends

.subckt nmos_1p2$$47342636_3v512x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.2772p pd=2.14u as=0.2772p ps=2.14u w=0.63u l=0.28u
.ends

.subckt ypredec1_3v512x8m81 ly[5] ly[4] ly[7] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_3v512x8m81_1/alatch_3v512x8m81_0/a
+ ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/a ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S
+ ly[3] M1_NWELL13_3v512x8m81_0/VSUBS pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ ypredec1_bot_3v512x8m81_0/alatch_3v512x8m81_0/a ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D
Xypredec1_xax8_3v512x8m81_0 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_0/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_5/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_1/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_6/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_2/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_3/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_4/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_xax8_3v512x8m81
Xypredec1_ys_3v512x8m81_0 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_0/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[3] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[3] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xpmos_1p2$$47109164_3v512x8m81_0 pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb nmos_5p04310591302056_3v512x8m81_1/D
+ pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S nmos_5p04310591302056_3v512x8m81_1/D
+ pmos_1p2$$47109164_3v512x8m81
Xypredec1_ys_3v512x8m81_1 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_6/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[4] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[4] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_2 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_2/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[5] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[5] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_bot_3v512x8m81_0 ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/alatch_3v512x8m81_0/a ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ ypredec1_bot_3v512x8m81
Xypredec1_ys_3v512x8m81_3 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[6] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[6] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_bot_3v512x8m81_1 ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/alatch_3v512x8m81_0/a ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ ypredec1_bot_3v512x8m81
Xypredec1_ys_3v512x8m81_4 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_5/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[0] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[0] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_bot_3v512x8m81_2 ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_1/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/a ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/S
+ ypredec1_bot_3v512x8m81_0/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_0/pmos_5p0431059130204_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb
+ ypredec1_bot_3v512x8m81_2/pmos_1p2$$46887980_3v512x8m81_1/pmos_5p0431059130204_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ ypredec1_bot_3v512x8m81
Xypredec1_ys_3v512x8m81_5 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_1/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[1] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[1] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_6 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_4/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[2] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[2] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_7 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_2/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[5] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[5] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_8 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_7/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[6] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[6] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_9 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_3/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[7] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[7] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xnmos_5p04310591302056_3v512x8m81_0 M1_NWELL13_3v512x8m81_0/VSUBS clk nmos_5p04310591302056_3v512x8m81_1/D
+ M1_NWELL13_3v512x8m81_0/VSUBS nmos_5p04310591302056_3v512x8m81
Xypredec1_ys_3v512x8m81_10 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_1/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[1] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[1] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xnmos_5p04310591302056_3v512x8m81_1 nmos_5p04310591302056_3v512x8m81_1/D men M1_NWELL13_3v512x8m81_0/VSUBS
+ M1_NWELL13_3v512x8m81_0/VSUBS nmos_5p04310591302056_3v512x8m81
Xypredec1_ys_3v512x8m81_11 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_4/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[2] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[2] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_12 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_0/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[3] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[3] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_13 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_6/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[4] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[4] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_14 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_5/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ry[0] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ry[0] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xypredec1_ys_3v512x8m81_15 ypredec1_xax8_3v512x8m81_0/ypredec1_xa_3v512x8m81_3/pmos_1p2$$47820844_3v512x8m81_2/pmos_5p04310591302061_3v512x8m81_0/D
+ M1_NWELL13_3v512x8m81_0/VSUBS ly[7] M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS
+ ly[7] ypredec1_ys_3v512x8m81_9/pmos_5p04310591302055_3v512x8m81_3/D M1_NWELL13_3v512x8m81_0/VSUBS
+ ypredec1_ys_3v512x8m81
Xnmos_1p2$$47342636_3v512x8m81_0 nmos_5p04310591302056_3v512x8m81_1/D ypredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb
+ M1_NWELL13_3v512x8m81_0/VSUBS M1_NWELL13_3v512x8m81_0/VSUBS nmos_1p2$$47342636_3v512x8m81
X0 a_5490_186# clk nmos_5p04310591302056_3v512x8m81_1/D pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S pfet_03v3 ad=0.1917p pd=1.425u as=0.34345p ps=1.71u w=1.065u l=0.28u
X1 nmos_5p04310591302056_3v512x8m81_1/D clk a_5176_186# pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S pfet_03v3 ad=0.34345p pd=1.71u as=0.19435p ps=1.43u w=1.065u l=0.28u
X2 a_5176_186# men pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S pfet_03v3 ad=0.19435p pd=1.43u as=0.59108p ps=3.24u w=1.065u l=0.28u
X3 pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S men a_5490_186# pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/S pfet_03v3 ad=0.59108p pd=3.24u as=0.1917p ps=1.425u w=1.065u l=0.28u
.ends

.subckt pmos_5p04310591302064_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.6322p pd=17.39u as=3.6322p ps=17.39u w=8.255u l=0.28u
.ends

.subckt pmos_1p2$$47503404_3v512x8m81 pmos_5p04310591302064_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302064_3v512x8m81_0/D w_n133_n65#
Xpmos_5p04310591302064_3v512x8m81_0 pmos_5p04310591302064_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302064_3v512x8m81_0/S pmos_5p04310591302064_3v512x8m81
.ends

.subckt nmos_5p04310591302066_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.4454p pd=7.45u as=1.4454p ps=7.45u w=3.285u l=0.28u
.ends

.subckt pmos_5p04310591302063_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.7016p pd=13.16u as=2.7016p ps=13.16u w=6.14u l=0.28u
.ends

.subckt pmos_1p2$$47504428_3v512x8m81 pmos_5p04310591302063_3v512x8m81_0/S a_n14_n34#
+ w_n133_n66# pmos_5p04310591302063_3v512x8m81_0/D
Xpmos_5p04310591302063_3v512x8m81_0 pmos_5p04310591302063_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302063_3v512x8m81_0/S pmos_5p04310591302063_3v512x8m81
.ends

.subckt nmos_5p04310591302065_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.0714p pd=5.75u as=1.0714p ps=5.75u w=2.435u l=0.28u
.ends

.subckt nmos_1p2$$47502380_3v512x8m81 nmos_5p04310591302065_3v512x8m81_0/S a_n14_n34#
+ nmos_5p04310591302065_3v512x8m81_0/D VSUBS
Xnmos_5p04310591302065_3v512x8m81_0 nmos_5p04310591302065_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302065_3v512x8m81_0/S VSUBS nmos_5p04310591302065_3v512x8m81
.ends

.subckt xpredec0_bot_3v512x8m81 nmos_5p04310591302066_3v512x8m81_0/D m1_n74_3354#
+ alatch_3v512x8m81_0/a m1_n74_3071# m1_n74_3213# nmos_1p2$$47502380_3v512x8m81_0/nmos_5p04310591302065_3v512x8m81_0/S
+ pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D alatch_3v512x8m81_0/vss
+ pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/S m1_n74_2930#
+ m2_800_2096# alatch_3v512x8m81_0/enb pmos_1p2$$47503404_3v512x8m81_0/pmos_5p04310591302064_3v512x8m81_0/S
+ alatch_3v512x8m81_0/vdd
Xpmos_1p2$$47503404_3v512x8m81_0 pmos_1p2$$47503404_3v512x8m81_0/pmos_5p04310591302064_3v512x8m81_0/S
+ alatch_3v512x8m81_0/ab nmos_5p04310591302066_3v512x8m81_0/D pmos_1p2$$47503404_3v512x8m81_0/pmos_5p04310591302064_3v512x8m81_0/S
+ pmos_1p2$$47503404_3v512x8m81
Xnmos_5p04310591302066_3v512x8m81_0 nmos_5p04310591302066_3v512x8m81_0/D alatch_3v512x8m81_0/ab
+ alatch_3v512x8m81_0/vss alatch_3v512x8m81_0/vss nmos_5p04310591302066_3v512x8m81
Xpmos_1p2$$47504428_3v512x8m81_0 pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/S
+ nmos_5p04310591302066_3v512x8m81_0/D pmos_1p2$$47503404_3v512x8m81_0/pmos_5p04310591302064_3v512x8m81_0/S
+ pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D pmos_1p2$$47504428_3v512x8m81
Xnmos_1p2$$47502380_3v512x8m81_0 nmos_1p2$$47502380_3v512x8m81_0/nmos_5p04310591302065_3v512x8m81_0/S
+ nmos_5p04310591302066_3v512x8m81_0/D pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ alatch_3v512x8m81_0/vss nmos_1p2$$47502380_3v512x8m81
Xalatch_3v512x8m81_0 alatch_3v512x8m81_0/enb alatch_3v512x8m81_0/en alatch_3v512x8m81_0/ab
+ alatch_3v512x8m81_0/a alatch_3v512x8m81_0/vss m2_800_2096# alatch_3v512x8m81_0/vdd
+ alatch_3v512x8m81
.ends

.subckt nmos_1p2$$46563372_3v512x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_1p2$$47641644_3v512x8m81 nmos_5p04310591302057_3v512x8m81_0/S nmos_5p04310591302057_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v512x8m81_0 nmos_5p04310591302057_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v512x8m81_0/S VSUBS nmos_5p04310591302057_3v512x8m81
.ends

.subckt pmos_5p04310591302067_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.1196p pd=15.06u as=3.1196p ps=15.06u w=7.09u l=0.28u
.ends

.subckt pmos_1p2$$47642668_3v512x8m81 pmos_5p04310591302067_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302067_3v512x8m81_0/D w_n194_n66#
Xpmos_5p04310591302067_3v512x8m81_0 pmos_5p04310591302067_3v512x8m81_0/D a_n14_n34#
+ w_n194_n66# pmos_5p04310591302067_3v512x8m81_0/S pmos_5p04310591302067_3v512x8m81
.ends

.subckt pmos_5p04310591302068_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt pmos_1p2$$47513644_3v512x8m81 pmos_5p04310591302068_3v512x8m81_0/S pmos_5p04310591302068_3v512x8m81_0/D
+ a_n14_n34# w_n133_n65#
Xpmos_5p04310591302068_3v512x8m81_0 pmos_5p04310591302068_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302068_3v512x8m81_0/S pmos_5p04310591302068_3v512x8m81
.ends

.subckt pmos_1p2$$47643692_3v512x8m81 w_n133_n66# pmos_5p04310591302067_3v512x8m81_0/S
+ a_n14_n34# pmos_5p04310591302067_3v512x8m81_0/D
Xpmos_5p04310591302067_3v512x8m81_0 pmos_5p04310591302067_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302067_3v512x8m81_0/S pmos_5p04310591302067_3v512x8m81
.ends

.subckt xpredec0_xa_3v512x8m81 m3_107_5938# m1_255_3759# a_612_1974# m1_255_3263#
+ m1_255_3619# m1_255_3901# pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D
+ m3_598_2319# a_472_3898# M3_M2$$47644716_3v512x8m81_2/VSUBS pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/S
+ nmos_1p2$$47641644_3v512x8m81_3/nmos_5p04310591302057_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D
+ nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
Xnmos_1p2$$47641644_3v512x8m81_0 nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ M3_M2$$47644716_3v512x8m81_2/VSUBS nmos_1p2$$47641644_3v512x8m81
Xpmos_1p2$$47642668_3v512x8m81_0 pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D
+ a_612_1974# pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47642668_3v512x8m81
Xnmos_1p2$$47641644_3v512x8m81_1 nmos_1p2$$47641644_3v512x8m81_3/nmos_5p04310591302057_3v512x8m81_0/D
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ M3_M2$$47644716_3v512x8m81_2/VSUBS nmos_1p2$$47641644_3v512x8m81
Xnmos_1p2$$47641644_3v512x8m81_2 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D
+ nmos_1p2$$47641644_3v512x8m81_3/nmos_5p04310591302057_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ M3_M2$$47644716_3v512x8m81_2/VSUBS nmos_1p2$$47641644_3v512x8m81
Xnmos_1p2$$47641644_3v512x8m81_3 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D
+ nmos_1p2$$47641644_3v512x8m81_3/nmos_5p04310591302057_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ M3_M2$$47644716_3v512x8m81_2/VSUBS nmos_1p2$$47641644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_0 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_1 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_2 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_3 pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_3/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47643692_3v512x8m81_0 pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S a_472_3898#
+ pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/D pmos_1p2$$47643692_3v512x8m81
X0 M3_M2$$47644716_3v512x8m81_2/VSUBS a_612_1974# a_539_2025# M3_M2$$47644716_3v512x8m81_2/VSUBS nfet_03v3 ad=3.1746p pd=12.55u as=1.0439p ps=6.085u w=5.72u l=0.28u
X1 a_539_2025# a_472_3898# pmos_1p2$$47643692_3v512x8m81_0/pmos_5p04310591302067_3v512x8m81_0/S M3_M2$$47644716_3v512x8m81_2/VSUBS nfet_03v3 ad=1.0439p pd=6.085u as=3.146p ps=12.54u w=5.72u l=0.28u
.ends

.subckt pmos_5p04310591302069_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt xpredec0_3v512x8m81 A[0] men x[0] x[1] x[2] clk xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ A[1] x[3] vdd vss xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
Xxpredec0_bot_3v512x8m81_0 xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D A[0] xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss vdd xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ a_4073_6932# pmos_5p04310591302069_3v512x8m81_0/D vdd vdd xpredec0_bot_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_0 a_4073_6932# pmos_5p04310591302069_3v512x8m81_0/D
+ vss vss nmos_1p2$$46563372_3v512x8m81
Xxpredec0_bot_3v512x8m81_1 xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D A[1] xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss vdd xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ a_4073_6932# pmos_5p04310591302069_3v512x8m81_0/D vdd vdd xpredec0_bot_3v512x8m81
Xxpredec0_xa_3v512x8m81_0 vss xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D
+ x[0] vdd xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss vdd vss vdd xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_xa_3v512x8m81
Xpmos_5p04310591302069_3v512x8m81_0 pmos_5p04310591302069_3v512x8m81_0/D a_4073_6932#
+ a_4073_6932# vdd vdd pmos_5p04310591302069_3v512x8m81
Xxpredec0_xa_3v512x8m81_2 vss xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D
+ x[1] vdd xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ vss vdd vss vdd xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_xa_3v512x8m81
Xxpredec0_xa_3v512x8m81_1 vss xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D
+ x[2] vdd xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D vss vdd
+ vss vdd xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_xa_3v512x8m81
Xxpredec0_xa_3v512x8m81_3 vss xpredec0_bot_3v512x8m81_1/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_0/pmos_1p2$$47504428_3v512x8m81_0/pmos_5p04310591302063_3v512x8m81_0/D
+ xpredec0_bot_3v512x8m81_0/nmos_5p04310591302066_3v512x8m81_0/D xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D
+ x[3] vdd xpredec0_bot_3v512x8m81_1/nmos_5p04310591302066_3v512x8m81_0/D vss vdd
+ vss vdd xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_xa_3v512x8m81
X0 vdd men a_3416_6773# vdd pfet_03v3 ad=0.448p pd=2.72u as=0.162p ps=1.205u w=0.8u l=0.28u
X1 vss clk a_4073_6932# vss nfet_03v3 ad=0.2794p pd=2.15u as=0.1651p ps=1.155u w=0.635u l=0.28u
X2 a_4073_6932# men vss vss nfet_03v3 ad=0.1651p pd=1.155u as=0.2794p ps=2.15u w=0.635u l=0.28u
X3 a_4073_6932# clk a_3091_6773# vdd pfet_03v3 ad=0.218p pd=1.345u as=0.208p ps=1.32u w=0.8u l=0.28u
X4 a_3091_6773# men vdd vdd pfet_03v3 ad=0.208p pd=1.32u as=0.364p ps=2.51u w=0.8u l=0.28u
X5 a_3416_6773# clk a_4073_6932# vdd pfet_03v3 ad=0.162p pd=1.205u as=0.218p ps=1.345u w=0.8u l=0.28u
.ends

.subckt pmos_5p04310591302072_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.1406p pd=10.61u as=2.1406p ps=10.61u w=4.865u l=0.28u
.ends

.subckt pmos_1p2$$47512620_3v512x8m81 pmos_5p04310591302072_3v512x8m81_0/D w_n133_n66#
+ a_n14_n34# pmos_5p04310591302072_3v512x8m81_0/S
Xpmos_5p04310591302072_3v512x8m81_0 pmos_5p04310591302072_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302072_3v512x8m81_0/S pmos_5p04310591302072_3v512x8m81
.ends

.subckt xpredec1_xa_3v512x8m81 m1_n40_n4147# m1_n40_n4005# m3_n46_n5510# a_145_n5643#
+ m1_n40_n3864# pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D
+ m1_n40_n3582# m1_n40_n3723# a_0_56# m1_n40_n3441# M2_M1$$47515692_3v512x8m81_3/VSUBS
+ a_465_n5643# pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S
+ a_305_n5643#
Xnmos_1p2$$47514668_3v512x8m81_0 M2_M1$$47515692_3v512x8m81_3/VSUBS pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D
+ pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S M2_M1$$47515692_3v512x8m81_3/VSUBS
+ nmos_1p2$$47514668_3v512x8m81
Xnmos_1p2$$47514668_3v512x8m81_1 pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D
+ M2_M1$$47515692_3v512x8m81_3/VSUBS pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ M2_M1$$47515692_3v512x8m81_3/VSUBS nmos_1p2$$47514668_3v512x8m81
Xnmos_1p2$$47514668_3v512x8m81_2 M2_M1$$47515692_3v512x8m81_3/VSUBS pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D
+ pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S M2_M1$$47515692_3v512x8m81_3/VSUBS
+ nmos_1p2$$47514668_3v512x8m81
Xpmos_1p2$$47512620_3v512x8m81_0 pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S a_145_n5643#
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47512620_3v512x8m81
Xpmos_1p2$$47512620_3v512x8m81_1 pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S a_465_n5643#
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47512620_3v512x8m81
Xpmos_1p2$$47512620_3v512x8m81_3 pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S a_305_n5643#
+ pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S pmos_1p2$$47512620_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_0 pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_1 pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47513644_3v512x8m81
Xpmos_1p2$$47513644_3v512x8m81_2 pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/D pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S
+ pmos_1p2$$47513644_3v512x8m81_2/pmos_5p04310591302068_3v512x8m81_0/S pmos_1p2$$47513644_3v512x8m81
X0 a_361_n5592# a_305_n5643# a_201_n5592# M2_M1$$47515692_3v512x8m81_3/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=1.5145p ps=6.345u w=5.825u l=0.28u
X1 a_201_n5592# a_145_n5643# M2_M1$$47515692_3v512x8m81_3/VSUBS M2_M1$$47515692_3v512x8m81_3/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=2.65037p ps=12.56u w=5.825u l=0.28u
X2 pmos_1p2$$47512620_3v512x8m81_3/pmos_5p04310591302072_3v512x8m81_0/S a_465_n5643# a_361_n5592# M2_M1$$47515692_3v512x8m81_3/VSUBS nfet_03v3 ad=2.82512p pd=12.62u as=1.5145p ps=6.345u w=5.825u l=0.28u
.ends

.subckt pmos_5p04310591302070_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.3528p pd=16.12u as=3.3528p ps=16.12u w=7.62u l=0.28u
.ends

.subckt pmos_1p2$$47337516_3v512x8m81 pmos_5p04310591302070_3v512x8m81_0/S pmos_5p04310591302070_3v512x8m81_0/D
+ a_n14_n34# w_n133_n65#
Xpmos_5p04310591302070_3v512x8m81_0 pmos_5p04310591302070_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302070_3v512x8m81_0/S pmos_5p04310591302070_3v512x8m81
.ends

.subckt nmos_5p04310591302071_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.3508p pd=7.02u as=1.3508p ps=7.02u w=3.07u l=0.28u
.ends

.subckt nmos_1p2$$47336492_3v512x8m81 nmos_5p04310591302071_3v512x8m81_0/S a_n14_n34#
+ nmos_5p04310591302071_3v512x8m81_0/D VSUBS
Xnmos_5p04310591302071_3v512x8m81_0 nmos_5p04310591302071_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302071_3v512x8m81_0/S VSUBS nmos_5p04310591302071_3v512x8m81
.ends

.subckt xpredec1_bot_3v512x8m81 m1_n74_2740# alatch_3v512x8m81_0/a pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D m1_n74_3446#
+ alatch_3v512x8m81_0/enb m1_n74_3164# m2_800_1786# alatch_3v512x8m81_0/vdd m1_n74_3305#
+ m1_n74_3023# alatch_3v512x8m81_0/vss m1_n74_2881# pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/S
Xpmos_1p2$$47337516_3v512x8m81_0 pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/S
+ pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/S pmos_1p2$$47337516_3v512x8m81
Xpmos_1p2$$47337516_3v512x8m81_1 pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/S
+ pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D alatch_3v512x8m81_0/ab
+ pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/S pmos_1p2$$47337516_3v512x8m81
Xnmos_1p2$$47336492_3v512x8m81_0 alatch_3v512x8m81_0/vss pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D alatch_3v512x8m81_0/vss
+ nmos_1p2$$47336492_3v512x8m81
Xnmos_1p2$$47336492_3v512x8m81_1 alatch_3v512x8m81_0/vss alatch_3v512x8m81_0/ab pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ alatch_3v512x8m81_0/vss nmos_1p2$$47336492_3v512x8m81
Xalatch_3v512x8m81_0 alatch_3v512x8m81_0/enb alatch_3v512x8m81_0/en alatch_3v512x8m81_0/ab
+ alatch_3v512x8m81_0/a alatch_3v512x8m81_0/vss m2_800_1786# alatch_3v512x8m81_0/vdd
+ alatch_3v512x8m81
.ends

.subckt xpredec1_3v512x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1]
+ A[0] clk w_5024_6624# xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd vdd vss
+ pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86# xpredec1_xa_3v512x8m81_7/m3_n46_n5510#
Xpmos_1p2$$47109164_3v512x8m81_0 pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb nmos_5p04310591302056_3v512x8m81_1/D
+ vdd nmos_5p04310591302056_3v512x8m81_1/D pmos_1p2$$47109164_3v512x8m81
Xxpredec1_xa_3v512x8m81_0 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[3] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_xa_3v512x8m81_1 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[1] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_xa_3v512x8m81_3 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[7] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_xa_3v512x8m81_2 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[5] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_bot_3v512x8m81_0 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ A[0] xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81
Xxpredec1_xa_3v512x8m81_4 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[2] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_bot_3v512x8m81_1 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ A[2] xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81
Xxpredec1_xa_3v512x8m81_5 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[0] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xxpredec1_bot_3v512x8m81_2 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ A[1] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ nmos_5p04310591302056_3v512x8m81_1/D xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81
Xnmos_5p04310591302056_3v512x8m81_0 vss clk nmos_5p04310591302056_3v512x8m81_1/D vss
+ nmos_5p04310591302056_3v512x8m81
Xxpredec1_xa_3v512x8m81_6 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[4] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xnmos_5p04310591302056_3v512x8m81_1 nmos_5p04310591302056_3v512x8m81_1/D men vss vss
+ nmos_5p04310591302056_3v512x8m81
Xxpredec1_xa_3v512x8m81_7 xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81_7/m3_n46_n5510# xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_0/pmos_5p04310591302070_3v512x8m81_0/D
+ x[6] xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_bot_3v512x8m81_0/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vss xpredec1_bot_3v512x8m81_1/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ vdd xpredec1_bot_3v512x8m81_2/pmos_1p2$$47337516_3v512x8m81_1/pmos_5p04310591302070_3v512x8m81_0/D
+ xpredec1_xa_3v512x8m81
Xnmos_1p2$$47342636_3v512x8m81_0 nmos_5p04310591302056_3v512x8m81_1/D xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/enb
+ vss vss nmos_1p2$$47342636_3v512x8m81
X0 a_5287_6723# men vdd w_5024_6624# pfet_03v3 ad=0.212p pd=1.46u as=0.5936p ps=3.24u w=1.06u l=0.28u
X1 a_5600_6723# clk nmos_5p04310591302056_3v512x8m81_1/D w_5024_6624# pfet_03v3 ad=0.19345p pd=1.425u as=0.32065p ps=1.665u w=1.06u l=0.28u
X2 nmos_5p04310591302056_3v512x8m81_1/D clk a_5287_6723# w_5024_6624# pfet_03v3 ad=0.32065p pd=1.665u as=0.212p ps=1.46u w=1.06u l=0.28u
X3 vdd men a_5600_6723# w_5024_6624# pfet_03v3 ad=0.5883p pd=3.23u as=0.19345p ps=1.425u w=1.06u l=0.28u
.ends

.subckt prexdec_top_3v512x8m81 A[2] xb[3] xa[0] xc[0] xc[1] xc[2] xc[3] xb[1] xb[2]
+ xb[0] xa[1] xa[2] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[1] xpredec0_3v512x8m81_1/xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec1_3v512x8m81_0/pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ xpredec1_3v512x8m81_0/clk xpredec0_3v512x8m81_1/xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_3v512x8m81_0/xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ A[4] A[5] xpredec0_3v512x8m81_0/xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ A[6] xpredec1_3v512x8m81_0/w_5024_6624# men xa[3] xpredec1_3v512x8m81_0/xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xpredec0_3v512x8m81_1/clk xpredec1_3v512x8m81_0/vdd VSUBS
Xxpredec0_3v512x8m81_0 A[3] men xb[0] xb[1] xb[2] xpredec0_3v512x8m81_1/clk xpredec0_3v512x8m81_0/xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ A[4] xb[3] xpredec1_3v512x8m81_0/vdd VSUBS xpredec0_3v512x8m81_0/xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_3v512x8m81
Xxpredec0_3v512x8m81_1 A[5] men xc[0] xc[1] xc[2] xpredec0_3v512x8m81_1/clk xpredec0_3v512x8m81_1/xpredec0_xa_3v512x8m81_2/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ A[6] xc[3] xpredec1_3v512x8m81_0/vdd VSUBS xpredec0_3v512x8m81_1/xpredec0_xa_3v512x8m81_3/nmos_1p2$$47641644_3v512x8m81_0/nmos_5p04310591302057_3v512x8m81_0/S
+ xpredec0_3v512x8m81
Xxpredec1_3v512x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] xpredec1_3v512x8m81_0/clk xpredec1_3v512x8m81_0/w_5024_6624# xpredec1_3v512x8m81_0/xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xpredec1_3v512x8m81_0/vdd VSUBS xpredec1_3v512x8m81_0/pmos_1p2$$47109164_3v512x8m81_0/pmos_5p04310591302062_3v512x8m81_0/w_n202_n86#
+ xpredec1_3v512x8m81_0/vdd xpredec1_3v512x8m81
.ends

.subckt nmos_5p04310591302090_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.465u
.ends

.subckt pmos_5p04310591302074_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.56u
.ends

.subckt nmos_5p04310591302085_3v512x8m81 a_530_n44# D a_n112_n44# a_209_n44# a_369_n44#
+ a_48_n44# S VSUBS
X0 D a_n112_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=2.0482p ps=10.19u w=4.655u l=0.28u
X1 S a_369_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=1.22192p ps=5.18u w=4.655u l=0.28u
X3 D a_530_n44# S VSUBS nfet_03v3 ad=2.0482p pd=10.19u as=1.22192p ps=5.18u w=4.655u l=0.28u
X4 S a_48_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
.ends

.subckt nmos_1p2$$48306220_3v512x8m81 nmos_5p04310591302085_3v512x8m81_0/S a_516_n34#
+ nmos_5p04310591302085_3v512x8m81_0/D a_195_n34# a_355_n34# a_n125_n34# a_34_n34#
+ VSUBS
Xnmos_5p04310591302085_3v512x8m81_0 a_516_n34# nmos_5p04310591302085_3v512x8m81_0/D
+ a_n125_n34# a_195_n34# a_355_n34# a_34_n34# nmos_5p04310591302085_3v512x8m81_0/S
+ VSUBS nmos_5p04310591302085_3v512x8m81
.ends

.subckt pmos_5p04310591302051_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6877p pd=3.165u as=1.1638p ps=6.17u w=2.645u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1638p pd=6.17u as=0.6877p ps=3.165u w=2.645u l=0.28u
.ends

.subckt pmos_5p04310591302094_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3872p pd=2.64u as=0.3872p ps=2.64u w=0.88u l=0.28u
.ends

.subckt pmos_1p2$$46285868_3v512x8m81 w_n133_n66# pmos_5p04310591302014_3v512x8m81_0/S
+ a_n14_n34# pmos_5p04310591302014_3v512x8m81_0/D
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt nmos_5p04310591302086_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6182p pd=3.69u as=0.6182p ps=3.69u w=1.405u l=0.28u
.ends

.subckt nmos_1p2$$48302124_3v512x8m81 nmos_5p04310591302086_3v512x8m81_0/S a_n14_n34#
+ nmos_5p04310591302086_3v512x8m81_0/D VSUBS
Xnmos_5p04310591302086_3v512x8m81_0 nmos_5p04310591302086_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302086_3v512x8m81_0/S VSUBS nmos_5p04310591302086_3v512x8m81
.ends

.subckt pmos_5p04310591302088_3v512x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=2.5608p ps=12.52u w=5.82u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=2.5608p pd=12.52u as=1.5132p ps=6.34u w=5.82u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
.ends

.subckt pmos_1p2$$202587180_3v512x8m81 pmos_5p04310591302014_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v512x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt pmos_5p04310591302079_3v512x8m81 D a_486_n44# a_165_n44# a_n156_n44# S a_4_n44#
+ a_646_n44# w_n330_n86# a_808_n44# a_325_n44#
X0 S a_646_n44# D w_n330_n86# pfet_03v3 ad=0.27162p pd=1.555u as=0.2665p ps=1.545u w=1.025u l=0.28u
X1 D a_165_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X2 D a_486_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X3 S a_4_n44# D w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X4 D a_n156_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.451p ps=2.93u w=1.025u l=0.28u
X5 S a_325_n44# D w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X6 D a_808_n44# S w_n330_n86# pfet_03v3 ad=0.451p pd=2.93u as=0.27162p ps=1.555u w=1.025u l=0.28u
.ends

.subckt nmos_5p04310591302039_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302020_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$202586156_3v512x8m81 pmos_5p04310591302014_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v512x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt nmos_1p2$$202595372_3v512x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt pmos_5p04310591302082_3v512x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X1 S a_662_n44# D w_n314_n86# pfet_03v3 ad=0.5082p pd=3.19u as=0.3003p ps=1.675u w=1.155u l=0.28u
X2 D a_502_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X3 S a_20_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X4 D a_181_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X5 D a_n140_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.5082p ps=3.19u w=1.155u l=0.28u
.ends

.subckt nmos_5p04310591302078_3v512x8m81 D S a_217_n44# a_n104_n44# a_56_n44# VSUBS
X0 D a_217_n44# S VSUBS nfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 S a_56_n44# D VSUBS nfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
X2 D a_n104_n44# S VSUBS nfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
.ends

.subckt nmos_1p2$$202596396_3v512x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302081_3v512x8m81 D a_634_n44# a_n168_n44# a_313_n44# a_795_n44#
+ a_474_n44# a_n8_n44# S a_153_n44# VSUBS
X0 D a_153_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X1 D a_474_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X2 D a_n168_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.28u
X3 S a_n8_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X4 D a_795_n44# S VSUBS nfet_03v3 ad=0.1826p pd=1.71u as=0.10892p ps=0.94u w=0.415u l=0.28u
X5 S a_313_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X6 S a_634_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
.ends

.subckt pmos_5p04310591302077_3v512x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.968p ps=5.28u w=2.2u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=0.968p pd=5.28u as=0.572p ps=2.72u w=2.2u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
.ends

.subckt nmos_5p04310591302075_3v512x8m81 D a_n252_n44# a_550_n44# a_229_n44# a_390_n44#
+ S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44# VSUBS
X0 D a_390_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X1 D a_n252_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.3938p ps=2.67u w=0.895u l=0.28u
X2 D a_69_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X3 S a_229_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X4 S a_550_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X5 S a_1192_n44# D VSUBS nfet_03v3 ad=0.3938p pd=2.67u as=0.2327p ps=1.415u w=0.895u l=0.28u
X6 D a_1032_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X7 S a_n92_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X8 S a_871_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X9 D a_711_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
.ends

.subckt pmos_5p04310591302080_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_5p04310591302076_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt wen_v2_3v512x8m81 IGWEN clk wen GWE vdd vss
Xpmos_1p2$$202587180_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_3/S pmos_5p04310591302014_3v512x8m81_4/D
+ pmos_5p04310591302041_3v512x8m81_1/S vdd pmos_1p2$$202587180_3v512x8m81
Xpmos_5p04310591302079_3v512x8m81_0 pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81_0/S vdd pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/S vdd pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302079_3v512x8m81
Xnmos_5p04310591302039_3v512x8m81_0 pmos_5p04310591302080_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_4/D
+ pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302041_3v512x8m81_0/S vss nmos_5p04310591302039_3v512x8m81
Xpmos_5p04310591302020_3v512x8m81_0 pmos_5p04310591302080_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_1/D
+ pmos_5p04310591302014_3v512x8m81_1/D vdd pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302020_3v512x8m81
Xpmos_1p2$$202586156_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_1/D pmos_5p04310591302014_3v512x8m81_2/S
+ vdd vdd pmos_1p2$$202586156_3v512x8m81
Xnmos_1p2$$202595372_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_1/S pmos_5p04310591302014_3v512x8m81_2/S
+ vss vss nmos_1p2$$202595372_3v512x8m81
Xnmos_1p2$$202595372_3v512x8m81_1 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302041_3v512x8m81_1/S
+ pmos_5p04310591302041_3v512x8m81_1/D vss nmos_1p2$$202595372_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_0 vdd pmos_5p04310591302079_3v512x8m81_0/D vdd pmos_5p04310591302041_3v512x8m81_0/D
+ pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302082_3v512x8m81_0 wen pmos_5p04310591302082_3v512x8m81_0/D wen wen
+ wen wen vdd wen vdd pmos_5p04310591302082_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_1 pmos_5p04310591302014_3v512x8m81_1/D clk vdd vdd
+ pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_2 vdd pmos_5p04310591302041_3v512x8m81_1/S vdd pmos_5p04310591302014_3v512x8m81_2/S
+ pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_3 vdd wen vdd pmos_5p04310591302014_3v512x8m81_3/S
+ pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_4 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302014_3v512x8m81_1/D
+ vdd vdd pmos_5p04310591302014_3v512x8m81
Xnmos_5p04310591302078_3v512x8m81_0 pmos_5p04310591302082_3v512x8m81_0/D vss wen wen
+ wen vss nmos_5p04310591302078_3v512x8m81
Xnmos_1p2$$202596396_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_2/S pmos_5p04310591302041_3v512x8m81_1/D
+ vss vss nmos_1p2$$202596396_3v512x8m81
Xpmos_5p04310591302041_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_4/D
+ vdd pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81
Xpmos_5p04310591302041_3v512x8m81_1 pmos_5p04310591302041_3v512x8m81_1/D pmos_5p04310591302014_3v512x8m81_1/D
+ vdd pmos_5p04310591302041_3v512x8m81_1/S pmos_5p04310591302041_3v512x8m81
Xnmos_5p04310591302081_3v512x8m81_0 pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81_0/S vss pmos_5p04310591302041_3v512x8m81_0/S
+ vss nmos_5p04310591302081_3v512x8m81
Xpmos_5p04310591302077_3v512x8m81_0 IGWEN pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302082_3v512x8m81_0/D vdd pmos_5p04310591302082_3v512x8m81_0/D vdd
+ pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302077_3v512x8m81
Xpmos_5p04310591302077_3v512x8m81_2 GWE pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302079_3v512x8m81_0/D vdd pmos_5p04310591302079_3v512x8m81_0/D vdd
+ pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302077_3v512x8m81
Xnmos_5p04310591302075_3v512x8m81_0 GWE pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D vss pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D
+ pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302079_3v512x8m81_0/D vss nmos_5p04310591302075_3v512x8m81
Xnmos_5p04310591302075_3v512x8m81_1 IGWEN pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D vss pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D
+ pmos_5p04310591302082_3v512x8m81_0/D pmos_5p04310591302082_3v512x8m81_0/D vss nmos_5p04310591302075_3v512x8m81
Xpmos_5p04310591302080_3v512x8m81_0 pmos_5p04310591302080_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_2/S
+ pmos_5p04310591302014_3v512x8m81_2/S vdd vdd pmos_5p04310591302080_3v512x8m81
Xnmos_5p04310591302010_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_1/S pmos_5p04310591302014_3v512x8m81_1/D
+ pmos_5p04310591302014_3v512x8m81_3/S vss nmos_5p04310591302010_3v512x8m81
Xnmos_5p04310591302076_3v512x8m81_0 pmos_5p04310591302080_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_2/S
+ pmos_5p04310591302014_3v512x8m81_2/S vss vss nmos_5p04310591302076_3v512x8m81
X0 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302014_3v512x8m81_1/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss wen pmos_5p04310591302014_3v512x8m81_3/S vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X2 pmos_5p04310591302014_3v512x8m81_1/D clk vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
X3 pmos_5p04310591302041_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_1/D pmos_5p04310591302041_3v512x8m81_0/S vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X4 vss pmos_5p04310591302079_3v512x8m81_0/D pmos_5p04310591302041_3v512x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt nmos_1p2$$48629804_3v512x8m81 nmos_5p04310591302039_3v512x8m81_0/S nmos_5p04310591302039_3v512x8m81_0/D
+ a_118_n34# a_n41_n34# VSUBS
Xnmos_5p04310591302039_3v512x8m81_0 nmos_5p04310591302039_3v512x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302039_3v512x8m81_0/S VSUBS nmos_5p04310591302039_3v512x8m81
.ends

.subckt pmos_5p04310591302087_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.6552p pd=22.04u as=4.6552p ps=22.04u w=10.58u l=0.28u
.ends

.subckt pmos_1p2$$47815724_3v512x8m81 pmos_5p04310591302087_3v512x8m81_0/D a_n14_n34#
+ pmos_5p04310591302087_3v512x8m81_0/S w_n133_n65#
Xpmos_5p04310591302087_3v512x8m81_0 pmos_5p04310591302087_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302087_3v512x8m81_0/S pmos_5p04310591302087_3v512x8m81
.ends

.subckt nmos_5p04310591302084_3v512x8m81 a_1394_n44# D a_2357_n44# a_1073_n44# a_2036_n44#
+ a_n51_n44# a_1715_n44# a_752_n44# a_n532_n44# a_431_n44# a_1554_n44# a_591_n44#
+ a_2197_n44# a_n211_n44# S a_110_n44# a_1876_n44# a_1233_n44# a_270_n44# a_912_n44#
+ a_2518_n44# a_n372_n44# VSUBS
X0 S a_270_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X1 D a_1715_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.90167p ps=3.96u w=3.435u l=0.28u
X2 D a_110_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X3 D a_2036_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X4 S a_n51_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X5 S a_591_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X6 D a_1073_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X7 D a_431_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X8 D a_2357_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X9 D a_1394_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X10 S a_n372_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X11 D a_752_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X12 S a_2518_n44# D VSUBS nfet_03v3 ad=1.5114p pd=7.75u as=0.90167p ps=3.96u w=3.435u l=0.28u
X13 S a_1233_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X14 S a_1876_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X15 D a_n211_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X16 S a_2197_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X17 S a_1554_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X18 D a_n532_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=1.5114p ps=7.75u w=3.435u l=0.28u
X19 S a_912_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
.ends

.subckt nmos_1p2$$48308268_3v512x8m81 nmos_5p04310591302084_3v512x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_2197_n44# nmos_5p04310591302084_3v512x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v512x8m81_0/D nmos_5p04310591302084_3v512x8m81_0/a_1233_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_1876_n44# nmos_5p04310591302084_3v512x8m81_0/a_n51_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_2518_n44# nmos_5p04310591302084_3v512x8m81_0/a_n372_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_752_n44# nmos_5p04310591302084_3v512x8m81_0/a_1394_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_2357_n44# nmos_5p04310591302084_3v512x8m81_0/a_431_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_591_n44# nmos_5p04310591302084_3v512x8m81_0/a_1073_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_2036_n44# nmos_5p04310591302084_3v512x8m81_0/S
+ nmos_5p04310591302084_3v512x8m81_0/a_110_n44# nmos_5p04310591302084_3v512x8m81_0/a_270_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_1715_n44# nmos_5p04310591302084_3v512x8m81_0/a_n532_n44#
+ VSUBS nmos_5p04310591302084_3v512x8m81_0/a_912_n44#
Xnmos_5p04310591302084_3v512x8m81_0 nmos_5p04310591302084_3v512x8m81_0/a_1394_n44#
+ nmos_5p04310591302084_3v512x8m81_0/D nmos_5p04310591302084_3v512x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_1073_n44# nmos_5p04310591302084_3v512x8m81_0/a_2036_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_n51_n44# nmos_5p04310591302084_3v512x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_752_n44# nmos_5p04310591302084_3v512x8m81_0/a_n532_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_431_n44# nmos_5p04310591302084_3v512x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_591_n44# nmos_5p04310591302084_3v512x8m81_0/a_2197_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_n211_n44# nmos_5p04310591302084_3v512x8m81_0/S
+ nmos_5p04310591302084_3v512x8m81_0/a_110_n44# nmos_5p04310591302084_3v512x8m81_0/a_1876_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_1233_n44# nmos_5p04310591302084_3v512x8m81_0/a_270_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_912_n44# nmos_5p04310591302084_3v512x8m81_0/a_2518_n44#
+ nmos_5p04310591302084_3v512x8m81_0/a_n372_n44# VSUBS nmos_5p04310591302084_3v512x8m81
.ends

.subckt nmos_5p04310591302093_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.56u
.ends

.subckt pmos_1p2$$47330348_3v512x8m81 pmos_5p04310591302041_3v512x8m81_0/D a_n14_89#
+ pmos_5p04310591302041_3v512x8m81_0/S w_n133_n65#
Xpmos_5p04310591302041_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81
.ends

.subckt pmos_5p04310591302089_3v512x8m81 a_2502_n44# a_1699_n44# D a_n67_n44# a_2341_n44#
+ a_1378_n44# a_2020_n44# a_1057_n44# a_n548_n44# a_94_n44# a_736_n44# a_n227_n44#
+ a_896_n44# w_n722_n86# S a_415_n44# a_2181_n44# a_1538_n44# a_575_n44# a_1860_n44#
+ a_1217_n44# a_n388_n44# a_254_n44#
X0 D a_n548_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=3.7708p ps=18.02u w=8.57u l=0.28u
X1 S a_575_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X2 D a_415_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X3 D a_1057_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X4 D a_2020_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X5 S a_896_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X6 D a_736_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X7 D a_1378_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X8 D a_2341_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X9 S a_n67_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X10 D a_1699_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.24962p ps=9.095u w=8.57u l=0.28u
X11 S a_2502_n44# D w_n722_n86# pfet_03v3 ad=3.7708p pd=18.02u as=2.24962p ps=9.095u w=8.57u l=0.28u
X12 S a_n388_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X13 S a_1217_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X14 S a_1860_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X15 S a_1538_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X16 S a_2181_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X17 D a_94_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X18 D a_n227_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X19 S a_254_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
.ends

.subckt pmos_5p04310591302073_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4563p pd=2.275u as=0.7722p ps=4.39u w=1.755u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7722p pd=4.39u as=0.4563p ps=2.275u w=1.755u l=0.28u
.ends

.subckt pmos_1p2$$48623660_3v512x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302073_3v512x8m81_0/D
+ a_118_n34# pmos_5p04310591302073_3v512x8m81_0/S
Xpmos_5p04310591302073_3v512x8m81_0 pmos_5p04310591302073_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302073_3v512x8m81_0/S pmos_5p04310591302073_3v512x8m81
.ends

.subckt pmos_5p04310591302092_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.465u
.ends

.subckt pmos_5p04310591302091_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.004p pd=19.08u as=4.004p ps=19.08u w=9.1u l=0.28u
.ends

.subckt pmos_1p2$$48624684_3v512x8m81 pmos_5p04310591302091_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302091_3v512x8m81_0/S
Xpmos_5p04310591302091_3v512x8m81_0 pmos_5p04310591302091_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302091_3v512x8m81_0/S pmos_5p04310591302091_3v512x8m81
.ends

.subckt pmos_5p0431059130203_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_1p2$$46273580_3v512x8m81 w_n133_n66# a_n42_n34# pmos_5p0431059130203_3v512x8m81_0/S
+ a_118_n34# pmos_5p0431059130203_3v512x8m81_0/D
Xpmos_5p0431059130203_3v512x8m81_0 pmos_5p0431059130203_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p0431059130203_3v512x8m81_0/S pmos_5p0431059130203_3v512x8m81
.ends

.subckt nmos_5p04310591302083_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1646p pd=1.64u as=0.1646p ps=1.64u w=0.35u l=0.28u
.ends

.subckt gen_3v512x8_3v512x8m81 VSS tblhl cen clk WEN GWE pmos_5p04310591302088_3v512x8m81_0/D
+ men IGWEN VDD wen_v2_3v512x8m81_0/wen
Xnmos_5p04310591302090_3v512x8m81_0 pmos_5p04310591302092_3v512x8m81_0/D pmos_5p04310591302074_3v512x8m81_1/D
+ VSS VSS nmos_5p04310591302090_3v512x8m81
Xpmos_5p04310591302074_3v512x8m81_0 pmos_5p04310591302074_3v512x8m81_0/D clk VDD VDD
+ pmos_5p04310591302074_3v512x8m81
Xpmos_5p04310591302074_3v512x8m81_1 pmos_5p04310591302074_3v512x8m81_1/D pmos_5p04310591302074_3v512x8m81_0/D
+ VDD VDD pmos_5p04310591302074_3v512x8m81
Xnmos_1p2$$48306220_3v512x8m81_0 VSS pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VSS nmos_1p2$$48306220_3v512x8m81
Xpmos_5p04310591302051_3v512x8m81_0 pmos_5p04310591302051_3v512x8m81_0/D pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S VDD VDD pmos_5p04310591302051_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_0 a_3546_5289# VSS pmos_1p2$$46285868_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ VSS nmos_1p2$$46563372_3v512x8m81
Xpmos_5p04310591302094_3v512x8m81_0 pmos_5p04310591302094_3v512x8m81_0/D pmos_5p04310591302092_3v512x8m81_0/D
+ VDD VDD pmos_5p04310591302094_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_1 pmos_5p04310591302051_3v512x8m81_0/D pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D
+ VSS VSS nmos_1p2$$46563372_3v512x8m81
Xpmos_1p2$$46285868_3v512x8m81_0 VDD VDD a_3546_5289# pmos_1p2$$46285868_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_1p2$$46285868_3v512x8m81
Xnmos_1p2$$46551084_3v512x8m81_0 pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ cen a_3546_5289# VSS nmos_1p2$$46551084_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_2 pmos_1p2$$46285868_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D
+ VSS nmos_1p2$$46563372_3v512x8m81
Xpmos_1p2$$46285868_3v512x8m81_1 VDD pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_1p2$$46285868_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D cen pmos_1p2$$46285868_3v512x8m81
Xnmos_1p2$$48302124_3v512x8m81_0 VSS pmos_5p04310591302094_3v512x8m81_0/D pmos_1p2$$48623660_3v512x8m81_0/pmos_5p04310591302073_3v512x8m81_0/D
+ VSS nmos_1p2$$48302124_3v512x8m81
Xpmos_5p04310591302088_3v512x8m81_0 pmos_5p04310591302088_3v512x8m81_0/D pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ VDD pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VDD pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_5p04310591302088_3v512x8m81
Xwen_v2_3v512x8m81_0 IGWEN clk wen_v2_3v512x8m81_0/wen GWE VDD VSS wen_v2_3v512x8m81
Xnmos_1p2$$48629804_3v512x8m81_0 VSS pmos_5p04310591302051_3v512x8m81_0/D pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S VSS nmos_1p2$$48629804_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_0 VDD tblhl pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S
+ VDD pmos_1p2$$47815724_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_1 pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VDD VDD pmos_1p2$$47815724_3v512x8m81
Xnmos_1p2$$48308268_3v512x8m81_0 pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D men pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D VSS pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D VSS pmos_5p04310591302088_3v512x8m81_0/D
+ nmos_1p2$$48308268_3v512x8m81
Xnmos_5p04310591302093_3v512x8m81_0 pmos_5p04310591302074_3v512x8m81_0/D clk VSS VSS
+ nmos_5p04310591302093_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_2 pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S
+ tblhl VDD VDD pmos_1p2$$47815724_3v512x8m81
Xnmos_5p04310591302093_3v512x8m81_1 pmos_5p04310591302074_3v512x8m81_1/D pmos_5p04310591302074_3v512x8m81_0/D
+ VSS VSS nmos_5p04310591302093_3v512x8m81
Xpmos_1p2$$47330348_3v512x8m81_0 pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D
+ a_3546_5289# pmos_1p2$$47330348_3v512x8m81_0/pmos_5p04310591302041_3v512x8m81_0/S
+ VDD pmos_1p2$$47330348_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_3 VDD pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S VDD pmos_1p2$$47815724_3v512x8m81
Xpmos_5p04310591302089_3v512x8m81_0 pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ men pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D VDD VDD pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302088_3v512x8m81_0/D
+ pmos_5p04310591302088_3v512x8m81_0/D pmos_5p04310591302089_3v512x8m81
Xpmos_1p2$$48623660_3v512x8m81_0 pmos_5p04310591302094_3v512x8m81_0/D VDD pmos_1p2$$48623660_3v512x8m81_0/pmos_5p04310591302073_3v512x8m81_0/D
+ pmos_5p04310591302094_3v512x8m81_0/D VDD pmos_1p2$$48623660_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_4 pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S VDD VDD pmos_1p2$$47815724_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_5 pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S VDD VDD pmos_1p2$$47815724_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_6 VDD pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VDD pmos_1p2$$47815724_3v512x8m81
Xpmos_1p2$$47815724_3v512x8m81_7 VDD pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S
+ pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VDD pmos_1p2$$47815724_3v512x8m81
Xnmos_1p2$$47342636_3v512x8m81_0 clk VSS a_3546_5289# VSS nmos_1p2$$47342636_3v512x8m81
Xpmos_5p04310591302092_3v512x8m81_0 pmos_5p04310591302092_3v512x8m81_0/D pmos_5p04310591302074_3v512x8m81_1/D
+ VDD VDD pmos_5p04310591302092_3v512x8m81
Xnmos_1p2$$47342636_3v512x8m81_1 men a_3546_5289# VSS VSS nmos_1p2$$47342636_3v512x8m81
Xpmos_1p2$$48624684_3v512x8m81_0 pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S
+ pmos_5p04310591302051_3v512x8m81_0/D VDD VDD pmos_1p2$$48624684_3v512x8m81
Xpmos_1p2$$48624684_3v512x8m81_1 pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S
+ pmos_1p2$$48623660_3v512x8m81_0/pmos_5p04310591302073_3v512x8m81_0/D VDD VDD pmos_1p2$$48624684_3v512x8m81
Xpmos_1p2$$46273580_3v512x8m81_0 VDD pmos_5p04310591302051_3v512x8m81_0/D VDD pmos_5p04310591302051_3v512x8m81_0/D
+ pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D pmos_1p2$$46273580_3v512x8m81
Xpmos_1p2$$48624684_3v512x8m81_2 VDD clk VDD pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S
+ pmos_1p2$$48624684_3v512x8m81
Xnmos_5p04310591302083_3v512x8m81_0 pmos_5p04310591302094_3v512x8m81_0/D pmos_5p04310591302092_3v512x8m81_0/D
+ VSS VSS nmos_5p04310591302083_3v512x8m81
X0 a_8790_2243# tblhl pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X1 a_3606_4291# men VDD VDD pfet_03v3 ad=0.2769p pd=1.585u as=0.50587p ps=3.08u w=1.065u l=0.28u
X2 a_7891_338# pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X3 a_6888_183# clk a_6728_183# VSS nfet_03v3 ad=2.7521p pd=11.105u as=2.7521p ps=11.105u w=10.585u l=0.28u
X4 VSS pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S a_7891_338# VSS nfet_03v3 ad=3.93622p pd=17.86u as=2.2009p ps=8.985u w=8.465u l=0.28u
X5 pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S tblhl a_8470_2243# VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X6 a_8470_2243# pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S VSS VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.96232p ps=5.14u w=2.115u l=0.28u
X7 pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S pmos_5p04310591302051_3v512x8m81_0/D a_6888_183# VSS nfet_03v3 ad=5.2925p pd=22.17u as=2.7521p ps=11.105u w=10.585u l=0.28u
X8 a_7571_338# pmos_1p2$$47815724_3v512x8m81_3/pmos_5p04310591302087_3v512x8m81_0/S VSS VSS nfet_03v3 ad=2.2009p pd=8.985u as=3.85157p ps=17.84u w=8.465u l=0.28u
X9 pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S pmos_1p2$$48624684_3v512x8m81_2/pmos_5p04310591302091_3v512x8m81_0/S a_7571_338# VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X10 a_6728_183# pmos_1p2$$48623660_3v512x8m81_0/pmos_5p04310591302073_3v512x8m81_0/D VSS VSS nfet_03v3 ad=2.7521p pd=11.105u as=4.6574p ps=22.05u w=10.585u l=0.28u
X11 a_3546_5289# clk a_3606_4291# VDD pfet_03v3 ad=0.50587p pd=3.08u as=0.2769p ps=1.585u w=1.065u l=0.28u
X12 VSS pmos_1p2$$47815724_3v512x8m81_7/pmos_5p04310591302087_3v512x8m81_0/S a_8790_2243# VSS nfet_03v3 ad=0.99405p pd=5.17u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt control_3v512x8_3v512x8m81 RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] A[0] CEN xb[1] xc[3] xc[1] xc[2]
+ xa[1] A[9] A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWEN ypredec1_3v512x8m81_0/ly[1]
+ ypredec1_3v512x8m81_0/ly[2] ypredec1_3v512x8m81_0/ly[4] ypredec1_3v512x8m81_0/ly[5]
+ ypredec1_3v512x8m81_0/ly[6] GWE ypredec1_3v512x8m81_0/ly[7] xa[0] prexdec_top_3v512x8m81_0/xpredec1_3v512x8m81_0/xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ xc[0] men VSS VDD
Xypredec1_3v512x8m81_0 ypredec1_3v512x8m81_0/ly[5] ypredec1_3v512x8m81_0/ly[4] ypredec1_3v512x8m81_0/ly[7]
+ ypredec1_3v512x8m81_0/ly[2] ypredec1_3v512x8m81_0/ly[1] LYS[7] RYS[0] RYS[1] RYS[2]
+ RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_3v512x8m81_0/ly[6] men A[0] A[1] A[2]
+ CLK A[2] A[1] VDD VDD VDD VDD VSS VDD A[0] VDD ypredec1_3v512x8m81
Xprexdec_top_3v512x8m81_0 A[5] xb[3] xa[0] xc[0] xc[1] xc[2] xc[3] xb[1] xb[2] xb[0]
+ xa[1] xa[2] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[4] VSS VDD CLK VSS VSS A[7] A[8]
+ VSS A[9] VDD men xa[3] prexdec_top_3v512x8m81_0/xpredec1_3v512x8m81_0/xpredec1_bot_3v512x8m81_2/alatch_3v512x8m81_0/vdd
+ CLK VDD VSS prexdec_top_3v512x8m81
Xgen_3v512x8_3v512x8m81_0 VSS tblhl CEN CLK gen_3v512x8_3v512x8m81_0/WEN GWE gen_3v512x8_3v512x8m81_0/pmos_5p04310591302088_3v512x8m81_0/D
+ men IGWEN VDD GWEN gen_3v512x8_3v512x8m81
.ends

.subckt x018SRAM_cell1_dummy_3v512x8m81 m3_82_330# a_248_342# a_248_592# w_82_512#
+ a_62_178# m2_346_89# m2_134_89# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_82_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_82_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt x018SRAM_cell1_cutPC_3v512x8m81 m3_82_330# a_248_342# a_248_592# a_62_178#
+ w_30_512# a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt array16_512_dummy_01_3v512x8m81 018SRAM_cell1_cutPC_3v512x8m81_34/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_53/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_14/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_30/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_53/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_19/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_63/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_24/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_42/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_24/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_63/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_15/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_0/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_49/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_44/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_11/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_44/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_44/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_54/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_54/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_40/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_15/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_29/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_25/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_25/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_32/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_25/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_4/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_48/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_35/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_21/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_54/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_37/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_52/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_16/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_55/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_16/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_50/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_26/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_26/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_35/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_31/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_46/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_56/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_17/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_56/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_17/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_1/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_16/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_27/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_27/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_45/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_12/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_37/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_37/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_41/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_47/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_57/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_18/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_61/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_1/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_18/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_26/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_59/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_28/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_28/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_45/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_22/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_1/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_38/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_51/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_19/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_58/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_19/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_36/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_29/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_29/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_36/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_43/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_49/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_40/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_17/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_49/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_59/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_59/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_46/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_42/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_3/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_27/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_6/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_47/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_10/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_23/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_56/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_2/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_20/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_20/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_53/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_30/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_30/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_40/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_42/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_50/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_35/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_7/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_21/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_60/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_21/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_62/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_5/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_18/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_31/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_3/a_62_178#
+ VSS VDD 018SRAM_cell1_cutPC_3v512x8m81_31/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_14/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_41/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_47/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_6/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_12/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_43/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_10/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_12/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_22/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_22/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_61/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_28/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_51/a_248_592#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_32/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_62/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_24/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_57/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_42/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_42/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_52/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_13/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_20/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_53/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_62/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_23/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_23/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_62/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_38/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_33/m3_82_330#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/a_248_342# 018SRAM_cell1_cutPC_3v512x8m81_50/a_248_592#
+ VSUBS 018SRAM_cell1_cutPC_3v512x8m81_43/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_34/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/a_248_592#
X018SRAM_cell1_cutPC_3v512x8m81_40 018SRAM_cell1_cutPC_3v512x8m81_40/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_40/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_40/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_51 018SRAM_cell1_cutPC_3v512x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_51/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_62 018SRAM_cell1_cutPC_3v512x8m81_62/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_62/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v512x8m81_62/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_62/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_30 018SRAM_cell1_cutPC_3v512x8m81_30/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_30/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_30/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_41 018SRAM_cell1_cutPC_3v512x8m81_41/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_41/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_41/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_52 018SRAM_cell1_cutPC_3v512x8m81_52/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_63 018SRAM_cell1_cutPC_3v512x8m81_63/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_63/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_42 018SRAM_cell1_cutPC_3v512x8m81_42/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_42/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_42/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_42/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_42/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_20 018SRAM_cell1_cutPC_3v512x8m81_20/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_20/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_42/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_20/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_42/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_53 018SRAM_cell1_cutPC_3v512x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_53/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_53/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_31 018SRAM_cell1_cutPC_3v512x8m81_31/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_31/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_32 018SRAM_cell1_cutPC_3v512x8m81_32/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_32/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_32/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_32/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_21 018SRAM_cell1_cutPC_3v512x8m81_21/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_21/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_21/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_41/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_43 018SRAM_cell1_cutPC_3v512x8m81_43/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_43/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_43/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_10 018SRAM_cell1_cutPC_3v512x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_10/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_54 018SRAM_cell1_cutPC_3v512x8m81_54/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_54/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_54/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_33 018SRAM_cell1_cutPC_3v512x8m81_33/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_33/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_33/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_22 018SRAM_cell1_cutPC_3v512x8m81_22/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_22/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_22/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_40/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_44 018SRAM_cell1_cutPC_3v512x8m81_44/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_44/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_44/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_11 018SRAM_cell1_cutPC_3v512x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_11/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_55 018SRAM_cell1_cutPC_3v512x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_34 018SRAM_cell1_cutPC_3v512x8m81_34/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_34/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_34/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_23 018SRAM_cell1_cutPC_3v512x8m81_23/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_23/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_23/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_45 018SRAM_cell1_cutPC_3v512x8m81_45/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_45/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_45/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_12 018SRAM_cell1_cutPC_3v512x8m81_12/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_12/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_12/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_56 018SRAM_cell1_cutPC_3v512x8m81_56/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_56/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_35 018SRAM_cell1_cutPC_3v512x8m81_35/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_35/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_35/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_24 018SRAM_cell1_cutPC_3v512x8m81_24/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_24/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_24/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_46 018SRAM_cell1_cutPC_3v512x8m81_46/m3_82_330# VSS
+ VDD 018SRAM_cell1_cutPC_3v512x8m81_46/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_13 018SRAM_cell1_cutPC_3v512x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_13/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_57 018SRAM_cell1_cutPC_3v512x8m81_57/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_57/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_36 018SRAM_cell1_cutPC_3v512x8m81_36/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_36/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_36/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_26 018SRAM_cell1_cutPC_3v512x8m81_26/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_26/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_26/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_36/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_37 018SRAM_cell1_cutPC_3v512x8m81_37/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_37/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_37/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_25 018SRAM_cell1_cutPC_3v512x8m81_25/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_25/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_25/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_37/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_47 018SRAM_cell1_cutPC_3v512x8m81_47/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_47/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_47/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_48 018SRAM_cell1_cutPC_3v512x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_48/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_15 018SRAM_cell1_cutPC_3v512x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_15/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_14 018SRAM_cell1_cutPC_3v512x8m81_14/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_14/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_58 018SRAM_cell1_cutPC_3v512x8m81_58/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_59 018SRAM_cell1_cutPC_3v512x8m81_59/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_59/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_27 018SRAM_cell1_cutPC_3v512x8m81_27/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_27/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_27/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_35/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_38 018SRAM_cell1_cutPC_3v512x8m81_38/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_38/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_38/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_38/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_16 018SRAM_cell1_cutPC_3v512x8m81_16/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_16/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_16/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_45/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_49 018SRAM_cell1_cutPC_3v512x8m81_49/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_49/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_49/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_28 018SRAM_cell1_cutPC_3v512x8m81_28/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_28/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_28/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_34/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_39 018SRAM_cell1_cutPC_3v512x8m81_39/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_39/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_39/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_39/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_17 018SRAM_cell1_cutPC_3v512x8m81_17/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_17/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_17/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_47/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_1 018SRAM_cell1_cutPC_3v512x8m81_1/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_1/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_1/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_1/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_29 018SRAM_cell1_cutPC_3v512x8m81_29/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_29/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_29/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_33/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_18 018SRAM_cell1_cutPC_3v512x8m81_18/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_18/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_18/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_44/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_0 018SRAM_cell1_cutPC_3v512x8m81_0/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_0/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v512x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_19 018SRAM_cell1_cutPC_3v512x8m81_19/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_19/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_19/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_43/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_2 018SRAM_cell1_cutPC_3v512x8m81_2/m3_82_330# VSS
+ 018SRAM_cell1_cutPC_3v512x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_2/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_3 018SRAM_cell1_cutPC_3v512x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_3/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_4 018SRAM_cell1_cutPC_3v512x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_5 018SRAM_cell1_cutPC_3v512x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_5/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_6 018SRAM_cell1_cutPC_3v512x8m81_6/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_7 018SRAM_cell1_cutPC_3v512x8m81_7/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_7/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_8 018SRAM_cell1_cutPC_3v512x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_9 018SRAM_cell1_cutPC_3v512x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_9/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_50 018SRAM_cell1_cutPC_3v512x8m81_50/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_50/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_50/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_60 018SRAM_cell1_cutPC_3v512x8m81_60/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
X018SRAM_cell1_cutPC_3v512x8m81_61 018SRAM_cell1_cutPC_3v512x8m81_61/m3_82_330# 018SRAM_cell1_cutPC_3v512x8m81_61/a_248_342#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v512x8m81_61/a_62_178#
+ 018SRAM_cell1_cutPC_3v512x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v512x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v512x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v512x8m81
.ends

.subckt new_dummyrow_unit_3v512x8m81 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
X018SRAM_cell1_dummy_3v512x8m81_6 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_7 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_8 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_9 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_10 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_11 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_12 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_13 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_14 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_15 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_1 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_0 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_2 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_3 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_4 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_5 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
.ends

.subckt new_dummyrowunit01_3v512x8m81 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# 018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89# 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89# VSUBS
X018SRAM_cell1_dummy_3v512x8m81_6 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_7 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_8 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_9 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_10 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_11 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_12 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_13 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_14 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_15 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_1 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_0 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_2 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_3 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_4 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_5 018SRAM_strap1_3v512x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
.ends

.subckt x018SRAM_cell1_3v512x8m81 m3_82_330# a_248_342# a_248_592# a_62_178# w_30_512#
+ a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt ldummy_3v512x4_3v512x8m81 array16_512_dummy_01_3v512x8m81_0/VSS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_17/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_17/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_46/m3_82_330#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/a_248_592#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_27/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_27/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_17/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_56/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_56/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_17/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_27/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_27/a_248_342#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/a_248_342#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_18/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_18/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/a_248_592# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/a_248_342#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_28/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_28/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_57/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_18/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_18/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_57/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_28/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_28/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/w_30_512#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/a_248_342#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_19/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/w_30_512# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_19/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/m3_82_330#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/a_248_342# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_29/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_58/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_19/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_58/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_19/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_29/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_29/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/w_30_512# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/w_30_512#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/w_30_512#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/a_248_592# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/m3_82_330# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/a_248_342# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_59/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_59/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_1/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/w_30_512# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_20/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_20/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_10/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_10/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_30/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_30/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_20/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_20/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_30/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/a_248_592#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_30/a_248_342#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/a_248_342#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_21/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_21/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_11/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_11/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_21/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_60/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_60/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_21/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/w_30_512# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_31/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_31/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/w_30_512#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/a_248_342# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_22/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_22/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_12/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_12/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_22/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_22/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/a_248_342#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_23/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_13/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_13/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_23/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_62/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_62/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_23/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/a_248_342#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_24/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_24/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_14/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_14/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_63/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_24/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_63/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_24/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/a_248_342# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_25/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_25/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_54/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_15/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_54/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_15/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_25/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_25/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_16/m2_346_89#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/a_248_342# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_16/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/m3_82_330# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/a_248_342# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_26/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_26/m2_134_89#
+ array16_512_dummy_01_3v512x8m81_0/VDD array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_55/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_16/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_16/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_55/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_26/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_26/a_248_342# 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/w_30_512# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/m3_82_330#
X018SRAM_cell1_dummy_3v512x8m81_6 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_7 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
Xarray16_512_dummy_01_3v512x8m81_0 VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/a_248_342#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_14/m3_82_330# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_14/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/a_248_342# VSUBS
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_63/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_24/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_24/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_63/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/a_248_592# VSUBS
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/a_248_342#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_54/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_15/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_54/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/a_248_342# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_15/a_248_342# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_8/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_25/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_25/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/w_30_512#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/w_30_512#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_55/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_16/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_55/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_16/a_248_342#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_26/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_26/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/m3_82_330#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/a_248_342#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/a_248_592#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_46/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/m3_82_330# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_56/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_0/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_17/m3_82_330#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_56/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_17/a_248_342# VSUBS
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_27/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_27/a_248_342# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_37/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/m3_82_330# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_9/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_1/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_57/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_57/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_18/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_1/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_18/a_248_342#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_28/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_28/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_45/w_30_512# VSUBS
+ VSUBS 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_38/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/m3_82_330# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_48/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_19/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_58/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_58/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_19/a_248_342# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_29/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_29/a_248_342#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_36/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/a_248_592# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/m3_82_330#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/a_248_592# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_59/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/a_248_342# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_59/a_248_342# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/a_248_592#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_10/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_47/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_10/a_248_342# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_2/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_20/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_20/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/w_30_512# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_4/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_30/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_30/m3_82_330#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_11/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_11/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_35/w_30_512#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_21/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_60/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_21/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_60/a_248_342# VSUBS
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_5/a_248_592# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_31/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/a_248_592#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/VSS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_31/a_248_342# 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/m3_82_330# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_41/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_12/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/a_248_342# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_12/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_22/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_22/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_61/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/w_30_512# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_6/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_51/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_32/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/w_30_512# array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_44/w_30_512# VSUBS
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_40/a_248_592# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_42/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_3/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_13/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_52/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_49/w_30_512# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_13/a_248_342#
+ VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_62/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_23/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_23/m3_82_330#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_62/a_248_342# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_53/w_30_512#
+ VSUBS array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_7/a_248_592#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_33/a_248_342#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_50/a_248_592# VSUBS
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_43/m3_82_330# array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_34/w_30_512#
+ array16_512_dummy_01_3v512x8m81_0/018SRAM_cell1_cutPC_3v512x8m81_39/a_248_592# array16_512_dummy_01_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_8 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_9 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
Xnew_dummyrow_unit_3v512x8m81_0 new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89#
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89# VSUBS
+ new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89# new_dummyrow_unit_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89#
+ VSUBS 018SRAM_cell1_3v512x8m81_1/w_30_512# new_dummyrow_unit_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_30 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_31 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_20 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_10 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_21 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_11 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_22 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_13 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_12 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_23 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_24 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_14 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_25 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_26 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_15 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_16 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_27 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_17 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_28 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_18 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_29 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_19 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
Xnew_dummyrowunit01_3v512x8m81_0 new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# VSUBS
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89# 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89#
+ new_dummyrowunit01_3v512x8m81_0/018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89# VSUBS
+ new_dummyrowunit01_3v512x8m81
X018SRAM_cell1_3v512x8m81_0 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD VSUBS
+ array16_512_dummy_01_3v512x8m81_0/VDD 018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_0 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_1 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_3v512x8m81_1 VSUBS VSUBS 018SRAM_cell1_3v512x8m81_1/w_30_512# VSUBS
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_2 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_3 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_4 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_5 VSUBS VSUBS array16_512_dummy_01_3v512x8m81_0/VDD
+ array16_512_dummy_01_3v512x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v512x8m81
.ends

.subckt dcap_103_novia_3v512x8m81 w_n205_0# a_n30_42# a_n119_86#
X0 a_n119_86# a_n30_42# a_n119_86# w_n205_0# pfet_03v3 ad=0.4717p pd=3.01u as=0 ps=0 w=1.06u l=1.74u
.ends

.subckt x018SRAM_cell1_2x_3v512x8m81 018SRAM_cell1_3v512x8m81_0/a_62_178# 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_3v512x8m81_1/a_62_178#
+ 018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_3v512x8m81_1/a_110_96#
X018SRAM_cell1_3v512x8m81_0 018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_3v512x8m81_0/a_62_178# 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_3v512x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v512x8m81
X018SRAM_cell1_3v512x8m81_1 018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_3v512x8m81_1/a_62_178# 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_3v512x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v512x8m81
.ends

.subckt Cell_array8x8_3v512x8m81 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178#
+ VSUBS
X018SRAM_cell1_2x_3v512x8m81_0[0|0] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|0] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|0] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|0] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|0] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|0] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|0] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|0] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|0] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|0] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|0] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|0] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|0] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|0] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|0] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|0] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|0] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|0] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|0] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|0] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|0] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|0] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|0] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|0] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|0] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|0] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|0] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|0] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|0] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|0] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|0] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|0] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|1] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|1] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|1] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|1] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|1] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|1] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|1] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|1] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|1] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|1] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|1] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|1] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|1] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|1] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|1] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|1] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|1] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|1] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|1] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|1] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|1] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|1] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|1] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|1] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|1] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|1] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|1] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|1] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|1] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|1] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|1] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|1] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|2] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|2] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|2] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|2] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|2] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|2] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|2] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|2] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|2] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|2] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|2] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|2] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|2] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|2] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|2] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|2] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|2] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|2] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|2] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|2] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|2] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|2] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|2] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|2] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|2] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|2] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|2] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|2] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|2] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|2] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|2] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|2] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|3] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|3] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|3] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|3] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|3] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|3] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|3] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|3] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|3] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|3] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|3] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|3] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|3] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|3] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|3] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|3] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|3] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|3] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|3] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|3] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|3] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|3] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|3] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|3] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|3] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|3] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|3] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|3] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|3] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|3] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|3] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|3] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|4] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|4] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|4] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|4] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|4] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|4] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|4] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|4] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|4] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|4] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|4] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|4] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|4] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|4] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|4] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|4] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|4] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|4] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|4] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|4] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|4] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|4] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|4] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|4] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|4] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|4] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|4] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|4] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|4] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|4] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|4] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|4] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|5] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|5] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|5] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|5] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|5] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|5] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|5] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|5] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|5] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|5] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|5] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|5] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|5] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|5] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|5] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|5] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|5] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|5] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|5] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|5] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|5] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|5] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|5] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|5] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|5] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|5] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|5] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|5] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|5] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|5] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|5] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|5] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|6] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|6] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|6] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|6] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|6] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|6] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|6] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|6] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|6] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|6] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|6] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|6] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|6] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|6] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|6] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|6] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|6] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|6] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|6] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|6] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|6] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|6] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|6] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|6] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|6] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|6] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|6] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|6] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|6] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|6] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|6] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|6] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[0|7] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[1|7] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[2|7] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[3|7] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[4|7] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[5|7] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[6|7] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[7|7] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[8|7] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[9|7] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[10|7] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[11|7] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[12|7] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[13|7] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[14|7] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[15|7] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[16|7] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[17|7] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[18|7] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[19|7] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[20|7] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[21|7] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[22|7] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[23|7] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[24|7] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[25|7] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[26|7] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[27|7] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[28|7] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[29|7] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[30|7] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0[31|7] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_0[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|0] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|0] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|0] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|0] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|0] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|0] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|0] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|0] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|0] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|0] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|0] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|0] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|0] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|0] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|0] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|0] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|0] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|0] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|0] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|0] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|0] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|0] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|0] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|0] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|0] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|0] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|0] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|0] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|0] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|0] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|0] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|0] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|1] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|1] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|1] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|1] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|1] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|1] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|1] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|1] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|1] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|1] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|1] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|1] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|1] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|1] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|1] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|1] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|1] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|1] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|1] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|1] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|1] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|1] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|1] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|1] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|1] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|1] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|1] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|1] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|1] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|1] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|1] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|1] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|2] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|2] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|2] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|2] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|2] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|2] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|2] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|2] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|2] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|2] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|2] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|2] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|2] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|2] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|2] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|2] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|2] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|2] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|2] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|2] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|2] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|2] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|2] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|2] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|2] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|2] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|2] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|2] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|2] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|2] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|2] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|2] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|3] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|3] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|3] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|3] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|3] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|3] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|3] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|3] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|3] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|3] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|3] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|3] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|3] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|3] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|3] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|3] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|3] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|3] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|3] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|3] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|3] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|3] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|3] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|3] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|3] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|3] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|3] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|3] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|3] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|3] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|3] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|3] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|4] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|4] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|4] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|4] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|4] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|4] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|4] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|4] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|4] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|4] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|4] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|4] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|4] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|4] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|4] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|4] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|4] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|4] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|4] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|4] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|4] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|4] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|4] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|4] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|4] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|4] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|4] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|4] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|4] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|4] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|4] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|4] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|5] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|5] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|5] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|5] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|5] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|5] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|5] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|5] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|5] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|5] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|5] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|5] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|5] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|5] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|5] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|5] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|5] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|5] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|5] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|5] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|5] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|5] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|5] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|5] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|5] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|5] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|5] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|5] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|5] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|5] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|5] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|5] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|6] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|6] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|6] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|6] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|6] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|6] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|6] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|6] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|6] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|6] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|6] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|6] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|6] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|6] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|6] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|6] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|6] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|6] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|6] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|6] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|6] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|6] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|6] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|6] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|6] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|6] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|6] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|6] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|6] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|6] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|6] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|6] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[0|7] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[1|7] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[2|7] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[3|7] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[4|7] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[5|7] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[6|7] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[7|7] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[8|7] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[9|7] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[10|7] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[11|7] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[12|7] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[13|7] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[14|7] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[15|7] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[16|7] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[17|7] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[18|7] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[19|7] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[20|7] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[21|7] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[22|7] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[23|7] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[24|7] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[25|7] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[26|7] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[27|7] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[28|7] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[29|7] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[30|7] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1[31|7] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_1[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|0] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|0] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|0] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|0] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|0] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|0] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|0] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|0] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|0] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|0] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|0] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|0] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|0] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|0] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|0] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|0] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|0] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|0] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|0] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|0] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|0] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|0] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|0] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|0] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|0] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|0] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|0] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|0] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|0] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|0] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|0] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|0] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|1] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|1] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|1] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|1] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|1] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|1] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|1] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|1] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|1] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|1] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|1] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|1] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|1] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|1] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|1] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|1] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|1] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|1] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|1] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|1] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|1] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|1] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|1] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|1] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|1] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|1] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|1] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|1] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|1] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|1] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|1] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|1] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|2] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|2] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|2] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|2] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|2] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|2] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|2] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|2] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|2] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|2] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|2] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|2] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|2] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|2] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|2] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|2] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|2] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|2] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|2] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|2] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|2] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|2] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|2] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|2] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|2] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|2] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|2] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|2] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|2] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|2] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|2] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|2] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|3] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|3] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|3] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|3] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|3] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|3] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|3] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|3] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|3] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|3] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|3] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|3] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|3] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|3] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|3] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|3] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|3] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|3] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|3] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|3] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|3] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|3] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|3] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|3] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|3] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|3] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|3] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|3] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|3] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|3] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|3] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|3] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|4] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|4] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|4] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|4] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|4] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|4] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|4] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|4] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|4] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|4] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|4] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|4] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|4] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|4] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|4] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|4] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|4] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|4] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|4] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|4] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|4] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|4] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|4] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|4] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|4] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|4] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|4] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|4] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|4] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|4] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|4] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|4] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|5] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|5] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|5] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|5] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|5] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|5] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|5] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|5] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|5] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|5] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|5] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|5] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|5] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|5] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|5] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|5] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|5] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|5] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|5] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|5] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|5] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|5] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|5] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|5] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|5] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|5] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|5] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|5] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|5] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|5] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|5] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|5] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|6] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|6] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|6] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|6] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|6] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|6] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|6] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|6] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|6] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|6] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|6] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|6] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|6] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|6] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|6] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|6] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|6] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|6] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|6] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|6] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|6] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|6] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|6] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|6] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|6] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|6] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|6] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|6] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|6] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|6] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|6] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|6] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[0|7] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[1|7] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[2|7] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[3|7] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[4|7] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[5|7] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[6|7] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[7|7] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[8|7] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[9|7] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[10|7] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[11|7] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[12|7] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[13|7] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[14|7] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[15|7] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[16|7] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[17|7] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[18|7] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[19|7] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[20|7] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[21|7] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[22|7] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[23|7] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[24|7] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[25|7] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[26|7] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[27|7] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[28|7] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[29|7] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[30|7] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2[31|7] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_2[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|0] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|0] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|0] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|0] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|0] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|0] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|0] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|0] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|0] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|0] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|0] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|0] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|0] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|0] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|0] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|0] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|0] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|0] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|0] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|0] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|0] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|0] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|0] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|0] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|0] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|0] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|0] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|0] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|0] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|0] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|0] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|0] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|0]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|1] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|1] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|1] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|1] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|1] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|1] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|1] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|1] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|1] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|1] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|1] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|1] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|1] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|1] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|1] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|1] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|1] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|1] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|1] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|1] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|1] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|1] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|1] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|1] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|1] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|1] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|1] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|1] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|1] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|1] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|1] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|1] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|1]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|2] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|2] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|2] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|2] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|2] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|2] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|2] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|2] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|2] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|2] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|2] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|2] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|2] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|2] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|2] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|2] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|2] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|2] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|2] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|2] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|2] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|2] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|2] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|2] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|2] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|2] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|2] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|2] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|2] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|2] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|2] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|2] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|2]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|3] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|3] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|3] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|3] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|3] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|3] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|3] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|3] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|3] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|3] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|3] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|3] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|3] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|3] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|3] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|3] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|3] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|3] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|3] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|3] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|3] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|3] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|3] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|3] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|3] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|3] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|3] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|3] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|3] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|3] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|3] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|3] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|3]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|4] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|4] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|4] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|4] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|4] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|4] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|4] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|4] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|4] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|4] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|4] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|4] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|4] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|4] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|4] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|4] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|4] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|4] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|4] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|4] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|4] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|4] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|4] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|4] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|4] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|4] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|4] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|4] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|4] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|4] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|4] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|4] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|4]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|5] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|5] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|5] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|5] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|5] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|5] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|5] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|5] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|5] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|5] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|5] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|5] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|5] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|5] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|5] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|5] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|5] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|5] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|5] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|5] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|5] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|5] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|5] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|5] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|5] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|5] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|5] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|5] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|5] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|5] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|5] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|5] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|5]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|6] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|6] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|6] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|6] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|6] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|6] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|6] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|6] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|6] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|6] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|6] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|6] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|6] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|6] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|6] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|6] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|6] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|6] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|6] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|6] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|6] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|6] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|6] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|6] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|6] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|6] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|6] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|6] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|6] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|6] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|6] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|6] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|6]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[0|7] 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[0]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[1|7] 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[1]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[2|7] 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[2]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[3|7] 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[3]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[4|7] 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[4]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[5|7] 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[5]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[6|7] 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[6]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[7|7] 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[7]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[8|7] 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[8]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[9|7] 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[10|7] 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[10]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[11|7] 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[11]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[12|7] 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[12]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[13|7] 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[13]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[14|7] 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[14]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[15|7] 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[15]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[16|7] 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[16]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[17|7] 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[17]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[18|7] 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[18]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[19|7] 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[19]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[20|7] 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[20]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[21|7] 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[21]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[22|7] 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[22]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[23|7] 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[23]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[24|7] 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[24]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[25|7] 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[25]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[26|7] 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[26]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[27|7] 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[27]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[28|7] 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[28]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[29|7] 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[29]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[30|7] 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[30]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3[31|7] 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v512x8m81_3[31]/018SRAM_strap1_3v512x8m81_1/a_91_178# 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v512x8m81_3[9]/018SRAM_strap1_3v512x8m81_1/w_91_512# 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ VSUBS 018SRAM_cell1_2x_3v512x8m81_3[9|7]/018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
.ends

.subckt nmos_5p04310591302011_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt pmos_5p0431059130206_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt pmos_1p2$$46885932_3v512x8m81 pmos_5p0431059130206_3v512x8m81_0/S pmos_5p0431059130206_3v512x8m81_0/D
+ a_118_89# a_n42_89# w_n133_n65#
Xpmos_5p0431059130206_3v512x8m81_0 pmos_5p0431059130206_3v512x8m81_0/D a_n42_89# a_118_89#
+ w_n133_n65# pmos_5p0431059130206_3v512x8m81_0/S pmos_5p0431059130206_3v512x8m81
.ends

.subckt pmos_5p0431059130209_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_5p0431059130207_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt nmos_1p2$$46884908_3v512x8m81 nmos_5p0431059130207_3v512x8m81_0/S a_n14_n34#
+ VSUBS nmos_5p0431059130207_3v512x8m81_0/D
Xnmos_5p0431059130207_3v512x8m81_0 nmos_5p0431059130207_3v512x8m81_0/D a_n14_n34#
+ nmos_5p0431059130207_3v512x8m81_0/S VSUBS nmos_5p0431059130207_3v512x8m81
.ends

.subckt pmos_5p0431059130201_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt pmos_1p2$$46889004_3v512x8m81 pmos_5p0431059130201_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v512x8m81_0/S
Xpmos_5p0431059130201_3v512x8m81_0 pmos_5p0431059130201_3v512x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v512x8m81_0/S pmos_5p0431059130201_3v512x8m81
.ends

.subckt nmos_5p0431059130205_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_1p2$$46883884_3v512x8m81 nmos_5p0431059130205_3v512x8m81_0/S nmos_5p0431059130205_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p0431059130205_3v512x8m81_0 nmos_5p0431059130205_3v512x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v512x8m81_0/S VSUBS nmos_5p0431059130205_3v512x8m81
.ends

.subckt din_3v512x8m81 d db datain wep men vdd vss pmos_5p0431059130206_3v512x8m81_0/D
+ m1_114_5647#
Xnmos_5p04310591302011_3v512x8m81_0 vss datain pmos_5p0431059130206_3v512x8m81_0/S
+ pmos_5p0431059130206_3v512x8m81_0/S vss nmos_5p04310591302011_3v512x8m81
Xnmos_5p04310591302011_3v512x8m81_1 nmos_5p04310591302011_3v512x8m81_1/D pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D
+ men pmos_5p0431059130206_3v512x8m81_0/S vss nmos_5p04310591302011_3v512x8m81
Xpmos_1p2$$46885932_3v512x8m81_0 pmos_5p0431059130206_3v512x8m81_0/S nmos_5p04310591302011_3v512x8m81_1/D
+ pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D men pmos_5p0431059130206_3v512x8m81_0/D
+ pmos_1p2$$46885932_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_0 pmos_5p0431059130201_3v512x8m81_0/S vss pmos_5p0431059130206_3v512x8m81_0/S
+ vss nmos_1p2$$46563372_3v512x8m81
Xnmos_1p2$$46563372_3v512x8m81_1 men vss pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D
+ vss nmos_1p2$$46563372_3v512x8m81
Xpmos_1p2$$46887980_3v512x8m81_0 vdd vdd pmos_5p0431059130201_3v512x8m81_0/S pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ pmos_1p2$$46887980_3v512x8m81
Xpmos_5p0431059130209_3v512x8m81_0 vdd pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ vdd pmos_5p0431059130209_3v512x8m81_0/S pmos_5p0431059130209_3v512x8m81
Xnmos_1p2$$46884908_3v512x8m81_0 vss pmos_5p0431059130201_3v512x8m81_0/S vss pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ nmos_1p2$$46884908_3v512x8m81
Xpmos_1p2$$46889004_3v512x8m81_0 pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ a_357_4344# vdd d pmos_1p2$$46889004_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_0 pmos_5p0431059130206_3v512x8m81_0/D nmos_5p04310591302011_3v512x8m81_1/D
+ pmos_5p0431059130206_3v512x8m81_0/D pmos_5p0431059130201_3v512x8m81_0/S pmos_5p0431059130201_3v512x8m81
Xnmos_1p2$$46883884_3v512x8m81_0 db pmos_5p0431059130209_3v512x8m81_0/S wep vss nmos_1p2$$46883884_3v512x8m81
Xpmos_1p2$$46889004_3v512x8m81_1 pmos_5p0431059130209_3v512x8m81_0/S a_357_4344# vdd
+ db pmos_1p2$$46889004_3v512x8m81
Xpmos_5p0431059130206_3v512x8m81_0 pmos_5p0431059130206_3v512x8m81_0/D datain pmos_5p0431059130206_3v512x8m81_0/S
+ pmos_5p0431059130206_3v512x8m81_0/D pmos_5p0431059130206_3v512x8m81_0/S pmos_5p0431059130206_3v512x8m81
Xnmos_1p2$$46883884_3v512x8m81_1 pmos_5p0431059130209_3v512x8m81_0/S vss pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ vss nmos_1p2$$46883884_3v512x8m81
Xnmos_5p04310591302010_3v512x8m81_0 vss nmos_5p04310591302011_3v512x8m81_1/D pmos_5p0431059130201_3v512x8m81_0/S
+ vss nmos_5p04310591302010_3v512x8m81
Xpmos_1p2$$46273580_3v512x8m81_0 pmos_5p0431059130206_3v512x8m81_0/D men pmos_5p0431059130206_3v512x8m81_0/D
+ men pmos_1p2$$46273580_3v512x8m81_0/pmos_5p0431059130203_3v512x8m81_0/D pmos_1p2$$46273580_3v512x8m81
Xnmos_1p2$$46883884_3v512x8m81_2 d pmos_1p2$$46889004_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ wep vss nmos_1p2$$46883884_3v512x8m81
Xpmos_1p2$$46273580_3v512x8m81_1 pmos_5p0431059130206_3v512x8m81_0/D pmos_5p0431059130201_3v512x8m81_0/S
+ pmos_5p0431059130206_3v512x8m81_0/D pmos_5p0431059130201_3v512x8m81_0/S pmos_5p0431059130206_3v512x8m81_0/S
+ pmos_1p2$$46273580_3v512x8m81
X0 vdd wep a_357_4344# vdd pfet_03v3 ad=0.38572p pd=2.5u as=0.1859p ps=1.23u w=0.695u l=0.28u
X1 a_357_4344# wep vdd vdd pfet_03v3 ad=0.1859p pd=1.23u as=0.38572p ps=2.5u w=0.695u l=0.28u
X2 a_357_4344# wep vss vss nfet_03v3 ad=0.28355p pd=2.13u as=0.3103p ps=2.23u w=0.535u l=0.28u
.ends

.subckt nmos_1p2$$202598444_3v512x8m81 nmos_5p04310591302010_3v512x8m81_0/S nmos_5p04310591302010_3v512x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302010_3v512x8m81_0 nmos_5p04310591302010_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v512x8m81_0/S VSUBS nmos_5p04310591302010_3v512x8m81
.ends

.subckt pmos_1p2$$202584108_3v512x8m81 pmos_5p04310591302014_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v512x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt nmos_5p04310591302042_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# VSUBS
X0 D a_265_n44# S VSUBS nfet_03v3 ad=0.1628p pd=1.62u as=97.125f ps=0.895u w=0.37u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=96.2f pd=0.89u as=0.1628p ps=1.62u w=0.37u l=0.28u
X2 S a_104_n44# D VSUBS nfet_03v3 ad=97.125f pd=0.895u as=96.2f ps=0.89u w=0.37u l=0.28u
.ends

.subckt nmos_1p2$$202594348_3v512x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
.ends

.subckt pmos_5p04310591302035_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$202583084_3v512x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302035_3v512x8m81_0/S
+ pmos_5p04310591302035_3v512x8m81_0/D a_118_n34#
Xpmos_5p04310591302035_3v512x8m81_0 pmos_5p04310591302035_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v512x8m81_0/S pmos_5p04310591302035_3v512x8m81
.ends

.subckt pmos_1p2$$202585132_3v512x8m81 pmos_5p04310591302014_3v512x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v512x8m81_0/D w_n119_n65#
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D a_n14_n34#
+ w_n119_n65# pmos_5p04310591302014_3v512x8m81_0/S pmos_5p04310591302014_3v512x8m81
.ends

.subckt pmos_5p04310591302043_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
.ends

.subckt wen_wm1_3v512x8m81 GWEN men wep wen vdd vss
Xnmos_1p2$$202598444_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_1/D pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302014_3v512x8m81_5/D vss nmos_1p2$$202598444_3v512x8m81
Xpmos_1p2$$202587180_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_1/D pmos_5p04310591302014_3v512x8m81_4/D
+ pmos_5p04310591302041_3v512x8m81_0/S vdd pmos_1p2$$202587180_3v512x8m81
Xnmos_5p04310591302039_3v512x8m81_0 men pmos_1p2$$202583084_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_1p2$$202583084_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D pmos_5p04310591302020_3v512x8m81_0/S
+ vss nmos_5p04310591302039_3v512x8m81
Xpmos_1p2$$202584108_3v512x8m81_0 pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/S vdd vdd pmos_1p2$$202584108_3v512x8m81
Xpmos_5p04310591302020_3v512x8m81_0 men pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D vdd pmos_5p04310591302020_3v512x8m81_0/S
+ pmos_5p04310591302020_3v512x8m81
Xpmos_1p2$$202586156_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_0/D pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ vdd vdd pmos_1p2$$202586156_3v512x8m81
Xnmos_1p2$$202595372_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302041_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/D vss nmos_1p2$$202595372_3v512x8m81
Xnmos_1p2$$202595372_3v512x8m81_1 pmos_5p04310591302041_3v512x8m81_0/S pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ vss vss nmos_1p2$$202595372_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_2/S wen vdd vdd
+ pmos_5p04310591302014_3v512x8m81
Xnmos_5p04310591302042_3v512x8m81_0 wep pmos_5p04310591302035_3v512x8m81_0/D vss pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_5p04310591302035_3v512x8m81_0/D vss nmos_5p04310591302042_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_1 pmos_5p04310591302014_3v512x8m81_1/D pmos_5p04310591302014_3v512x8m81_2/D
+ vdd vdd pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_2 pmos_5p04310591302014_3v512x8m81_2/D GWEN vdd
+ pmos_5p04310591302014_3v512x8m81_2/S pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_3 pmos_5p04310591302014_3v512x8m81_5/S men vdd vdd
+ pmos_5p04310591302014_3v512x8m81
Xnmos_1p2$$202594348_3v512x8m81_0 pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_1p2$$202583084_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D vss vss nmos_1p2$$202594348_3v512x8m81
Xpmos_1p2$$202583084_3v512x8m81_0 pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ vdd vdd pmos_1p2$$202583084_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_1p2$$202583084_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_4 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302014_3v512x8m81_5/D
+ vdd vdd pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_5 pmos_5p04310591302014_3v512x8m81_5/D vss vdd pmos_5p04310591302014_3v512x8m81_5/S
+ pmos_5p04310591302014_3v512x8m81
Xnmos_1p2$$202596396_3v512x8m81_0 pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ vss pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D vss nmos_1p2$$202596396_3v512x8m81
Xnmos_1p2$$202596396_3v512x8m81_1 pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ pmos_5p04310591302041_3v512x8m81_0/D vss vss nmos_1p2$$202596396_3v512x8m81
Xpmos_5p04310591302041_3v512x8m81_0 pmos_5p04310591302041_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_5/D
+ vdd pmos_5p04310591302041_3v512x8m81_0/S pmos_5p04310591302041_3v512x8m81
Xpmos_5p04310591302035_3v512x8m81_0 pmos_5p04310591302035_3v512x8m81_0/D pmos_5p04310591302020_3v512x8m81_0/S
+ pmos_5p04310591302020_3v512x8m81_0/S vdd vdd pmos_5p04310591302035_3v512x8m81
Xpmos_1p2$$202585132_3v512x8m81_0 vdd pmos_1p2$$202584108_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/S
+ pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D vdd pmos_1p2$$202585132_3v512x8m81
Xpmos_5p04310591302043_3v512x8m81_0 wep pmos_5p04310591302035_3v512x8m81_0/D vdd pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_5p04310591302035_3v512x8m81_0/D vdd pmos_5p04310591302043_3v512x8m81
Xnmos_5p04310591302010_3v512x8m81_0 vss pmos_1p2$$202585132_3v512x8m81_0/pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_5p04310591302020_3v512x8m81_0/S vss nmos_5p04310591302010_3v512x8m81
X0 pmos_5p04310591302014_3v512x8m81_5/D men vss vss nfet_03v3 ad=0.1651p pd=1.155u as=0.2794p ps=2.15u w=0.635u l=0.28u
X1 vss GWEN pmos_5p04310591302014_3v512x8m81_2/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
X2 pmos_5p04310591302014_3v512x8m81_4/D pmos_5p04310591302014_3v512x8m81_5/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X3 pmos_5p04310591302014_3v512x8m81_1/D pmos_5p04310591302014_3v512x8m81_2/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X4 vss vss pmos_5p04310591302014_3v512x8m81_5/D vss nfet_03v3 ad=0.2794p pd=2.15u as=0.1651p ps=1.155u w=0.635u l=0.28u
X5 pmos_5p04310591302035_3v512x8m81_0/D pmos_5p04310591302020_3v512x8m81_0/S vss vss nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
X6 pmos_5p04310591302014_3v512x8m81_2/D wen vss vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p0431059130200_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt nmos_1p2$$47119404_3v512x8m81 nmos_5p0431059130200_3v512x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v512x8m81_0/S VSUBS
Xnmos_5p0431059130200_3v512x8m81_0 nmos_5p0431059130200_3v512x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v512x8m81_0/S VSUBS nmos_5p0431059130200_3v512x8m81
.ends

.subckt nmos_5p0431059130202_3v512x8m81 D a_n32_n44# a_136_n44# S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=91.3f pd=0.92u as=0.1561p ps=1.64u w=0.265u l=0.28u
X1 S a_136_n44# D VSUBS nfet_03v3 ad=0.15742p pd=1.65u as=91.3f ps=0.92u w=0.265u l=0.28u
.ends

.subckt ypass_gate_a_3v512x8m81 vss b bb ypass pcb m3_n41_6881# a_64_7110# m3_n41_5924#
+ m3_n41_6639# m3_n41_4610# vdd pmos_5p0431059130201_3v512x8m81_0/D m3_n41_5682# via1_2_3v512x8m81_0/VSUBS
+ pmos_5p0431059130201_3v512x8m81_1/D pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ m3_n41_5198# m3_n41_5440# m3_n41_6156#
Xnmos_1p2$$47119404_3v512x8m81_1 pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass pmos_5p0431059130201_3v512x8m81_0/D via1_2_3v512x8m81_0/VSUBS nmos_1p2$$47119404_3v512x8m81
Xnmos_1p2$$47119404_3v512x8m81_3 pmos_5p0431059130201_3v512x8m81_1/D ypass bb via1_2_3v512x8m81_0/VSUBS
+ nmos_1p2$$47119404_3v512x8m81
Xnmos_5p0431059130202_3v512x8m81_0 nmos_5p0431059130202_3v512x8m81_0/D ypass ypass
+ via1_2_3v512x8m81_0/VSUBS via1_2_3v512x8m81_0/VSUBS nmos_5p0431059130202_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_0 pmos_5p0431059130201_3v512x8m81_0/D pcb vdd bb
+ pmos_5p0431059130201_3v512x8m81
Xpmos_1p2$$46889004_3v512x8m81_1 pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ nmos_5p0431059130202_3v512x8m81_0/D vdd pmos_5p0431059130201_3v512x8m81_0/D pmos_1p2$$46889004_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_1 pmos_5p0431059130201_3v512x8m81_1/D nmos_5p0431059130202_3v512x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v512x8m81
X0 vdd pcb pmos_5p0431059130201_3v512x8m81_0/D vdd pfet_03v3 ad=1.06988p pd=4.52u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 pmos_5p0431059130201_3v512x8m81_0/D pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.99855p ps=4.43u w=1.585u l=0.28u
X2 vdd ypass nmos_5p0431059130202_3v512x8m81_0/D vdd pfet_03v3 ad=0.5143p pd=2.87u as=0.34055p ps=1.675u w=0.695u l=0.28u
X3 vdd pcb bb vdd pfet_03v3 ad=1.07325p pd=4.53u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=1.0017p ps=4.44u w=1.59u l=0.28u
X5 nmos_5p0431059130202_3v512x8m81_0/D ypass vdd vdd pfet_03v3 ad=0.34055p pd=1.675u as=0.38572p ps=2.5u w=0.695u l=0.28u
.ends

.subckt ypass_gate_3v512x8m81 vss b bb ypass pcb m3_n41_6881# db m3_n41_5924# m3_n41_6639#
+ m3_n41_4610# vdd pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ m3_n41_5682# a_94_7110# m3_n41_5198# m3_n41_5440# m3_n41_6156# via1_2_3v512x8m81_0/VSUBS
Xnmos_1p2$$47119404_3v512x8m81_1 pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass b via1_2_3v512x8m81_0/VSUBS nmos_1p2$$47119404_3v512x8m81
Xnmos_1p2$$47119404_3v512x8m81_3 db ypass bb via1_2_3v512x8m81_0/VSUBS nmos_1p2$$47119404_3v512x8m81
Xnmos_5p0431059130202_3v512x8m81_0 nmos_5p0431059130202_3v512x8m81_0/D ypass ypass
+ via1_2_3v512x8m81_0/VSUBS via1_2_3v512x8m81_0/VSUBS nmos_5p0431059130202_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_0 b pcb vdd bb pmos_5p0431059130201_3v512x8m81
Xpmos_1p2$$46889004_3v512x8m81_1 pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ nmos_5p0431059130202_3v512x8m81_0/D vdd b pmos_1p2$$46889004_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_1 db nmos_5p0431059130202_3v512x8m81_0/D vdd bb pmos_5p0431059130201_3v512x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.92722p pd=4.34u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 b pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.93515p ps=4.35u w=1.585u l=0.28u
X2 nmos_5p0431059130202_3v512x8m81_0/D ypass vdd vdd pfet_03v3 ad=0.26235p pd=1.45u as=0.46218p ps=2.72u w=0.695u l=0.28u
X3 vdd ypass nmos_5p0431059130202_3v512x8m81_0/D vdd pfet_03v3 ad=0.39963p pd=2.54u as=0.26235p ps=1.45u w=0.695u l=0.28u
X4 vdd pcb bb vdd pfet_03v3 ad=0.93015p pd=4.35u as=0.4134p ps=2.11u w=1.59u l=0.28u
X5 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=0.9381p ps=4.36u w=1.59u l=0.28u
.ends

.subckt mux821_3v512x8m81 ypass_gate_3v512x8m81_1/bb ypass_gate_3v512x8m81_4/b ypass_gate_3v512x8m81_1/db
+ ypass_gate_3v512x8m81_2/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_5/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_6/b ypass_gate_a_3v512x8m81_0/ypass ypass_gate_3v512x8m81_6/bb
+ ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D ypass_gate_3v512x8m81_3/bb
+ ypass_gate_3v512x8m81_7/db ypass_gate_3v512x8m81_5/db ypass_gate_3v512x8m81_1/b
+ ypass_gate_3v512x8m81_3/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_a_3v512x8m81_0/bb ypass_gate_3v512x8m81_6/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_1/ypass ypass_gate_3v512x8m81_3/b ypass_gate_3v512x8m81_2/ypass
+ ypass_gate_3v512x8m81_3/ypass ypass_gate_3v512x8m81_5/b ypass_gate_3v512x8m81_4/ypass
+ ypass_gate_3v512x8m81_5/ypass ypass_gate_3v512x8m81_5/bb ypass_gate_3v512x8m81_2/bb
+ ypass_gate_3v512x8m81_4/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_6/ypass ypass_gate_3v512x8m81_7/b ypass_gate_3v512x8m81_7/ypass
+ ypass_gate_3v512x8m81_4/db ypass_gate_3v512x8m81_1/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_a_3v512x8m81_0/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_7/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_2/b ypass_gate_3v512x8m81_7/bb
+ ypass_gate_3v512x8m81_4/bb ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
Xypass_gate_a_3v512x8m81_0 ypass_gate_3v512x8m81_7/vss ypass_gate_a_3v512x8m81_0/b
+ ypass_gate_a_3v512x8m81_0/bb ypass_gate_a_3v512x8m81_0/ypass ypass_gate_3v512x8m81_7/pcb
+ ypass_gate_3v512x8m81_7/m3_n41_6881# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5924#
+ ypass_gate_3v512x8m81_7/m3_n41_6639# ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd
+ ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D ypass_gate_3v512x8m81_7/m3_n41_5682#
+ VSUBS ypass_gate_3v512x8m81_1/db ypass_gate_a_3v512x8m81_0/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5198# ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156#
+ ypass_gate_a_3v512x8m81
Xypass_gate_3v512x8m81_1 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_1/b ypass_gate_3v512x8m81_1/bb
+ ypass_gate_3v512x8m81_1/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_1/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_1/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_2 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_2/b ypass_gate_3v512x8m81_2/bb
+ ypass_gate_3v512x8m81_2/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_4/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_2/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_3 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_3/b ypass_gate_3v512x8m81_3/bb
+ ypass_gate_3v512x8m81_3/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_5/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_3/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_4 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_4/b ypass_gate_3v512x8m81_4/bb
+ ypass_gate_3v512x8m81_4/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_4/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_4/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_5 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_5/b ypass_gate_3v512x8m81_5/bb
+ ypass_gate_3v512x8m81_5/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_5/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_5/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_6 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_6/b ypass_gate_3v512x8m81_6/bb
+ ypass_gate_3v512x8m81_6/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_7/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_6/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
Xypass_gate_3v512x8m81_7 ypass_gate_3v512x8m81_7/vss ypass_gate_3v512x8m81_7/b ypass_gate_3v512x8m81_7/bb
+ ypass_gate_3v512x8m81_7/ypass ypass_gate_3v512x8m81_7/pcb ypass_gate_3v512x8m81_7/m3_n41_6881#
+ ypass_gate_3v512x8m81_7/db ypass_gate_3v512x8m81_7/m3_n41_5924# ypass_gate_3v512x8m81_7/m3_n41_6639#
+ ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/vdd ypass_gate_3v512x8m81_7/pmos_1p2$$46889004_3v512x8m81_1/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_7/m3_n41_5682# ypass_gate_3v512x8m81_7/a_94_7110# ypass_gate_3v512x8m81_7/m3_n41_5198#
+ ypass_gate_3v512x8m81_7/m3_n41_5440# ypass_gate_3v512x8m81_7/m3_n41_6156# VSUBS
+ ypass_gate_3v512x8m81
.ends

.subckt nmos_5p04310591302012_3v512x8m81 a_n83_n44# D a_77_n44# S a_237_n44# a_397_n44#
+ VSUBS
X0 S a_77_n44# D VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_397_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_237_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X3 D a_n83_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$45107244_3v512x8m81 a_223_n34# a_383_n34# nmos_5p04310591302012_3v512x8m81_0/S
+ a_n96_n34# a_63_n34# VSUBS nmos_5p04310591302012_3v512x8m81_0/D
Xnmos_5p04310591302012_3v512x8m81_0 a_n96_n34# nmos_5p04310591302012_3v512x8m81_0/D
+ a_63_n34# nmos_5p04310591302012_3v512x8m81_0/S a_223_n34# a_383_n34# VSUBS nmos_5p04310591302012_3v512x8m81
.ends

.subckt nmos_5p04310591302016_3v512x8m81 a_124_n45# a_284_n45# D a_446_n45# a_768_n45#
+ a_n198_n45# a_n38_n45# a_606_n45# S a_928_n45# VSUBS
X0 S a_928_n45# D VSUBS nfet_03v3 ad=0.7155p pd=4.08u as=0.4134p ps=2.11u w=1.59u l=0.28u
X1 D a_n198_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.70755p ps=4.07u w=1.59u l=0.28u
X2 S a_n38_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X3 S a_606_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 D a_768_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X5 D a_446_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X6 S a_284_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X7 D a_124_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46552108_3v512x8m81 nmos_5p04310591302016_3v512x8m81_0/D nmos_5p04310591302016_3v512x8m81_0/a_606_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_n198_n45# nmos_5p04310591302016_3v512x8m81_0/a_928_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_124_n45# nmos_5p04310591302016_3v512x8m81_0/a_284_n45#
+ nmos_5p04310591302016_3v512x8m81_0/S nmos_5p04310591302016_3v512x8m81_0/a_446_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_768_n45# nmos_5p04310591302016_3v512x8m81_0/a_n38_n45#
+ VSUBS
Xnmos_5p04310591302016_3v512x8m81_0 nmos_5p04310591302016_3v512x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_284_n45# nmos_5p04310591302016_3v512x8m81_0/D
+ nmos_5p04310591302016_3v512x8m81_0/a_446_n45# nmos_5p04310591302016_3v512x8m81_0/a_768_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_n198_n45# nmos_5p04310591302016_3v512x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v512x8m81_0/a_606_n45# nmos_5p04310591302016_3v512x8m81_0/S
+ nmos_5p04310591302016_3v512x8m81_0/a_928_n45# VSUBS nmos_5p04310591302016_3v512x8m81
.ends

.subckt pmos_5p04310591302019_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46898220_3v512x8m81 w_n133_n66# pmos_5p04310591302019_3v512x8m81_0/D
+ a_n14_84# pmos_5p04310591302019_3v512x8m81_0/S
Xpmos_5p04310591302019_3v512x8m81_0 pmos_5p04310591302019_3v512x8m81_0/D a_n14_84#
+ w_n133_n66# pmos_5p04310591302019_3v512x8m81_0/S pmos_5p04310591302019_3v512x8m81
.ends

.subckt nmos_5p04310591302017_3v512x8m81 a_n37_n44# D a_929_n44# a_125_n44# a_285_n44#
+ a_447_n44# a_769_n44# S a_607_n44# a_n197_n44# VSUBS
X0 D a_769_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X1 D a_447_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X2 D a_n197_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X3 S a_n37_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X4 S a_285_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X5 D a_125_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X6 S a_929_n44# D VSUBS nfet_03v3 ad=0.58963p pd=3.54u as=0.3445p ps=1.845u w=1.325u l=0.28u
X7 S a_607_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_1p2$$46550060_3v512x8m81 a_915_n34# nmos_5p04310591302017_3v512x8m81_0/D
+ a_111_n34# a_271_n34# a_433_n34# a_593_n34# a_n51_n34# a_755_n34# a_n210_n34# nmos_5p04310591302017_3v512x8m81_0/S
+ VSUBS
Xnmos_5p04310591302017_3v512x8m81_0 a_n51_n34# nmos_5p04310591302017_3v512x8m81_0/D
+ a_915_n34# a_111_n34# a_271_n34# a_433_n34# a_755_n34# nmos_5p04310591302017_3v512x8m81_0/S
+ a_593_n34# a_n210_n34# VSUBS nmos_5p04310591302017_3v512x8m81
.ends

.subckt pmos_5p04310591302013_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46286892_3v512x8m81 w_n133_n66# pmos_5p04310591302013_3v512x8m81_0/S
+ pmos_5p04310591302013_3v512x8m81_0/D a_n70_n34# a_90_n34# a_251_n34#
Xpmos_5p04310591302013_3v512x8m81_0 pmos_5p04310591302013_3v512x8m81_0/D a_251_n34#
+ pmos_5p04310591302013_3v512x8m81_0/S a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302013_3v512x8m81
.ends

.subckt pmos_5p04310591302018_3v512x8m81 a_20_n45# D a_181_n45# a_502_n45# a_662_n45#
+ a_n140_n45# S a_341_n45# w_n314_n86#
X0 S a_341_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_662_n45# D w_n314_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_502_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 S a_20_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_181_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X5 D a_n140_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46549036_3v512x8m81 a_327_n34# w_n188_n50# a_488_n34# a_n154_n34#
+ pmos_5p04310591302018_3v512x8m81_0/S a_167_n34# a_6_n34# pmos_5p04310591302018_3v512x8m81_0/D
+ a_648_n34#
Xpmos_5p04310591302018_3v512x8m81_0 a_6_n34# pmos_5p04310591302018_3v512x8m81_0/D
+ a_167_n34# a_488_n34# a_648_n34# a_n154_n34# pmos_5p04310591302018_3v512x8m81_0/S
+ a_327_n34# w_n188_n50# pmos_5p04310591302018_3v512x8m81
.ends

.subckt pmos_5p04310591302021_3v512x8m81 a_76_n44# D a_n84_n44# w_n258_n86# S a_237_n44#
+ a_397_n44#
X0 S a_397_n44# D w_n258_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1092p ps=0.94u w=0.42u l=0.28u
X1 D a_237_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.11025p ps=0.945u w=0.42u l=0.28u
X2 D a_n84_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.1848p ps=1.72u w=0.42u l=0.28u
X3 S a_76_n44# D w_n258_n86# pfet_03v3 ad=0.11025p pd=0.945u as=0.1092p ps=0.94u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46896172_3v512x8m81 w_n133_n66# pmos_5p04310591302021_3v512x8m81_0/a_237_n44#
+ pmos_5p04310591302021_3v512x8m81_0/a_397_n44# pmos_5p04310591302021_3v512x8m81_0/a_76_n44#
+ pmos_5p04310591302021_3v512x8m81_0/S pmos_5p04310591302021_3v512x8m81_0/D pmos_5p04310591302021_3v512x8m81_0/a_n84_n44#
Xpmos_5p04310591302021_3v512x8m81_0 pmos_5p04310591302021_3v512x8m81_0/a_76_n44# pmos_5p04310591302021_3v512x8m81_0/D
+ pmos_5p04310591302021_3v512x8m81_0/a_n84_n44# w_n133_n66# pmos_5p04310591302021_3v512x8m81_0/S
+ pmos_5p04310591302021_3v512x8m81_0/a_237_n44# pmos_5p04310591302021_3v512x8m81_0/a_397_n44#
+ pmos_5p04310591302021_3v512x8m81
.ends

.subckt pmos_1p2$$46897196_3v512x8m81 w_n133_n66# pmos_5p04310591302020_3v512x8m81_0/S
+ a_n42_n34# pmos_5p04310591302020_3v512x8m81_0/D a_118_n34#
Xpmos_5p04310591302020_3v512x8m81_0 pmos_5p04310591302020_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302020_3v512x8m81_0/S pmos_5p04310591302020_3v512x8m81
.ends

.subckt nmos_5p04310591302015_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6996p pd=4.06u as=0.6996p ps=4.06u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46553132_3v512x8m81 nmos_5p04310591302015_3v512x8m81_0/S a_n14_n34#
+ nmos_5p04310591302015_3v512x8m81_0/D VSUBS
Xnmos_5p04310591302015_3v512x8m81_0 nmos_5p04310591302015_3v512x8m81_0/D a_n14_n34#
+ nmos_5p04310591302015_3v512x8m81_0/S VSUBS nmos_5p04310591302015_3v512x8m81
.ends

.subckt sa_3v512x8m81 qp wep se pcb vdd vss d
Xnmos_1p2$$45107244_3v512x8m81_0 qp qp qp pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ qp vss vss nmos_1p2$$45107244_3v512x8m81
Xnmos_1p2$$46552108_3v512x8m81_0 nmos_1p2$$46552108_3v512x8m81_0/nmos_5p04310591302016_3v512x8m81_0/D
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S vss nmos_1p2$$46552108_3v512x8m81
Xpmos_1p2$$46898220_3v512x8m81_0 d pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ d d pmos_1p2$$46898220_3v512x8m81
Xnmos_1p2$$46550060_3v512x8m81_0 se nmos_1p2$$46552108_3v512x8m81_0/nmos_5p04310591302016_3v512x8m81_0/D
+ se se se se se se se vss vss nmos_1p2$$46550060_3v512x8m81
Xpmos_1p2$$46898220_3v512x8m81_1 d d d pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81
Xpmos_1p2$$46286892_3v512x8m81_0 d d d pcb pcb pcb pmos_1p2$$46286892_3v512x8m81
Xnmos_1p2$$46551084_3v512x8m81_0 qp vss pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ vss nmos_1p2$$46551084_3v512x8m81
Xpmos_1p2$$46285868_3v512x8m81_0 d pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pcb pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46285868_3v512x8m81
Xpmos_1p2$$46549036_3v512x8m81_0 qp vdd pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S vdd qp pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ qp pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46549036_3v512x8m81
Xpmos_1p2$$46896172_3v512x8m81_0 d pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S d pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ pmos_1p2$$46896172_3v512x8m81
Xpmos_1p2$$46897196_3v512x8m81_0 d d se pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ se pmos_1p2$$46897196_3v512x8m81
Xpmos_1p2$$46897196_3v512x8m81_1 d d se pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ se pmos_1p2$$46897196_3v512x8m81
Xpmos_1p2$$46897196_3v512x8m81_2 d d se pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ se pmos_1p2$$46897196_3v512x8m81
Xpmos_1p2$$46897196_3v512x8m81_3 d d se pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ se pmos_1p2$$46897196_3v512x8m81
Xnmos_1p2$$46553132_3v512x8m81_0 pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_3v512x8m81
Xnmos_1p2$$46553132_3v512x8m81_1 vss vss pmos_1p2$$46898220_3v512x8m81_1/pmos_5p04310591302019_3v512x8m81_0/S
+ vss nmos_1p2$$46553132_3v512x8m81
.ends

.subckt nmos_5p04310591302026_3v512x8m81 a_154_n44# D a_n168_n44# a_476_n44# a_798_n44#
+ a_314_n44# a_n8_n44# S a_636_n44# VSUBS
X0 S a_636_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_314_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_n168_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X3 S a_n8_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_798_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X5 D a_476_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X6 D a_154_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$45102124_3v512x8m81 a_140_n34# a_462_n34# nmos_5p04310591302026_3v512x8m81_0/S
+ a_n181_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v512x8m81_0/D a_622_n34#
+ a_n22_n34# VSUBS
Xnmos_5p04310591302026_3v512x8m81_0 a_140_n34# nmos_5p04310591302026_3v512x8m81_0/D
+ a_n181_n34# a_462_n34# a_784_n34# a_300_n34# a_n22_n34# nmos_5p04310591302026_3v512x8m81_0/S
+ a_622_n34# VSUBS nmos_5p04310591302026_3v512x8m81
.ends

.subckt pmos_1p2$$46284844_3v512x8m81 w_n133_n66# pmos_5p04310591302035_3v512x8m81_0/S
+ a_118_n34# pmos_5p04310591302035_3v512x8m81_0/D a_n42_n34#
Xpmos_5p04310591302035_3v512x8m81_0 pmos_5p04310591302035_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v512x8m81_0/S pmos_5p04310591302035_3v512x8m81
.ends

.subckt nmos_5p04310591302023_3v512x8m81 D a_n32_n44# a_136_n44# S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=92.8f pd=0.92u as=0.1576p ps=1.64u w=0.28u l=0.28u
X1 S a_136_n44# D VSUBS nfet_03v3 ad=0.159p pd=1.65u as=92.8f ps=0.92u w=0.28u l=0.28u
.ends

.subckt nmos_5p04310591302028_3v512x8m81 D a_64_n44# a_226_n44# a_386_n44# a_548_n44#
+ S a_n96_n44# VSUBS
X0 D a_548_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X1 S a_386_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_226_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X3 D a_n96_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X4 S a_64_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302025_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n85#
X0 D a_265_n44# S w_n230_n85# pfet_03v3 ad=0.9306p pd=5.11u as=0.55518p ps=2.64u w=2.115u l=0.28u
X1 D a_n56_n44# S w_n230_n85# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X2 S a_104_n44# D w_n230_n85# pfet_03v3 ad=0.55518p pd=2.64u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$46281772_3v512x8m81 w_n133_n66# pmos_5p04310591302025_3v512x8m81_0/S
+ a_251_n34# a_n70_n34# pmos_5p04310591302025_3v512x8m81_0/D a_90_n34#
Xpmos_5p04310591302025_3v512x8m81_0 pmos_5p04310591302025_3v512x8m81_0/D a_251_n34#
+ pmos_5p04310591302025_3v512x8m81_0/S a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302025_3v512x8m81
.ends

.subckt pmos_5p04310591302038_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.2464p pd=2u as=0.2464p ps=2u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302037_3v512x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X1 S a_662_n44# D VSUBS nfet_03v3 ad=0.5852p pd=3.54u as=0.3458p ps=1.85u w=1.33u l=0.28u
X2 D a_502_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X3 S a_20_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X4 D a_181_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X5 D a_n140_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.5852p ps=3.54u w=1.33u l=0.28u
.ends

.subckt nmos_1p2$$45103148_3v512x8m81 a_327_n34# a_n153_n34# a_488_n34# a_167_n34#
+ nmos_5p04310591302037_3v512x8m81_0/S a_6_n34# a_648_n34# nmos_5p04310591302037_3v512x8m81_0/D
+ VSUBS
Xnmos_5p04310591302037_3v512x8m81_0 a_6_n34# nmos_5p04310591302037_3v512x8m81_0/D
+ a_167_n34# a_488_n34# a_648_n34# a_n153_n34# nmos_5p04310591302037_3v512x8m81_0/S
+ a_327_n34# VSUBS nmos_5p04310591302037_3v512x8m81
.ends

.subckt pmos_5p04310591302030_3v512x8m81 a_871_n45# D a_n252_n45# a_550_n45# a_229_n45#
+ w_n426_n86# a_390_n45# S a_n92_n45# a_1032_n45# a_1192_n45# a_711_n45# a_69_n45#
X0 D a_390_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X1 D a_n252_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.5566p ps=3.41u w=1.265u l=0.28u
X2 D a_69_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X3 S a_229_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X4 S a_550_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X5 S a_1192_n45# D w_n426_n86# pfet_03v3 ad=0.5566p pd=3.41u as=0.3289p ps=1.785u w=1.265u l=0.28u
X6 D a_1032_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X7 S a_n92_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X8 S a_871_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X9 D a_711_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
.ends

.subckt pmos_1p2$$45095980_3v512x8m81 a_697_n34# a_n106_n34# a_n266_n34# a_376_n34#
+ pmos_5p04310591302030_3v512x8m81_0/D a_1018_n34# a_1178_n34# a_55_n34# w_987_n66#
+ a_857_n34# a_536_n34# pmos_5p04310591302030_3v512x8m81_0/S a_215_n34#
Xpmos_5p04310591302030_3v512x8m81_0 a_857_n34# pmos_5p04310591302030_3v512x8m81_0/D
+ a_n266_n34# a_536_n34# a_215_n34# w_987_n66# a_376_n34# pmos_5p04310591302030_3v512x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34# a_55_n34# pmos_5p04310591302030_3v512x8m81
.ends

.subckt pmos_5p04310591302027_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt pmos_5p04310591302024_3v512x8m81 w_n286_n86# a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S
X0 D a_n112_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_369_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_209_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 D a_530_n44# S w_n286_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X4 S a_48_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46282796_3v512x8m81 a_n126_n34# pmos_5p04310591302024_3v512x8m81_0/S
+ a_195_n34# a_516_n34# w_163_n66# pmos_5p04310591302024_3v512x8m81_0/D a_355_n34#
+ a_34_n34#
Xpmos_5p04310591302024_3v512x8m81_0 w_163_n66# a_516_n34# pmos_5p04310591302024_3v512x8m81_0/D
+ a_n126_n34# a_195_n34# a_355_n34# a_34_n34# pmos_5p04310591302024_3v512x8m81_0/S
+ pmos_5p04310591302024_3v512x8m81
.ends

.subckt nmos_5p04310591302029_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.54067p pd=3.32u as=0.3159p ps=1.735u w=1.215u l=0.28u
.ends

.subckt nmos_1p2$$45100076_3v512x8m81 nmos_5p04310591302029_3v512x8m81_0/S a_118_n34#
+ nmos_5p04310591302029_3v512x8m81_0/D a_n41_n34# VSUBS
Xnmos_5p04310591302029_3v512x8m81_0 nmos_5p04310591302029_3v512x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302029_3v512x8m81_0/S VSUBS nmos_5p04310591302029_3v512x8m81
.ends

.subckt nmos_5p04310591302032_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.23585p pd=1.95u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_5p04310591302022_3v512x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.8382p ps=4.69u w=1.905u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=0.8382p pd=4.69u as=0.4953p ps=2.425u w=1.905u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
.ends

.subckt pmos_1p2$$46283820_3v512x8m81 pmos_5p04310591302022_3v512x8m81_0/D a_536_n34#
+ a_215_n34# a_697_n34# a_n106_n34# a_n266_n34# a_376_n34# pmos_5p04310591302022_3v512x8m81_0/S
+ w_984_n66# a_1018_n34# a_1178_n34# a_55_n34# a_857_n34#
Xpmos_5p04310591302022_3v512x8m81_0 pmos_5p04310591302022_3v512x8m81_0/D a_n266_n34#
+ a_536_n34# a_215_n34# w_984_n66# a_376_n34# pmos_5p04310591302022_3v512x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34# a_55_n34# a_857_n34# pmos_5p04310591302022_3v512x8m81
.ends

.subckt nmos_5p04310591302036_3v512x8m81 a_530_n44# D a_n112_n44# a_209_n44# a_369_n44#
+ a_48_n44# S VSUBS
X0 D a_n112_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_369_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.13913p ps=1.055u w=0.53u l=0.28u
X3 D a_530_n44# S VSUBS nfet_03v3 ad=0.2332p pd=1.94u as=0.13913p ps=1.055u w=0.53u l=0.28u
X4 S a_48_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt nmos_1p2$$45101100_3v512x8m81 a_195_n34# a_35_n34# nmos_5p04310591302036_3v512x8m81_0/S
+ a_516_n34# a_n125_n34# nmos_5p04310591302036_3v512x8m81_0/D a_356_n34# VSUBS
Xnmos_5p04310591302036_3v512x8m81_0 a_516_n34# nmos_5p04310591302036_3v512x8m81_0/D
+ a_n125_n34# a_195_n34# a_356_n34# a_35_n34# nmos_5p04310591302036_3v512x8m81_0/S
+ VSUBS nmos_5p04310591302036_3v512x8m81
.ends

.subckt nmos_5p04310591302033_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.28u
.ends

.subckt pmos_5p04310591302031_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4134p pd=2.11u as=0.6996p ps=4.06u w=1.59u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6996p pd=4.06u as=0.4134p ps=2.11u w=1.59u l=0.28u
.ends

.subckt pmos_1p2$$46287916_3v512x8m81 w_n133_n66# a_n42_n34# pmos_5p04310591302031_3v512x8m81_0/S
+ pmos_5p04310591302031_3v512x8m81_0/D a_118_n34#
Xpmos_5p04310591302031_3v512x8m81_0 pmos_5p04310591302031_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302031_3v512x8m81_0/S pmos_5p04310591302031_3v512x8m81
.ends

.subckt sacntl_2_3v512x8m81 pcb se pmos_5p04310591302027_3v512x8m81_2/S pmos_5p04310591302027_3v512x8m81_1/S
+ men vdd vss
Xnmos_1p2$$45102124_3v512x8m81_0 pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S vss pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pcb pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ vss nmos_1p2$$45102124_3v512x8m81
Xpmos_1p2$$46284844_3v512x8m81_0 vdd vdd pmos_5p04310591302027_3v512x8m81_1/S pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_5p04310591302027_3v512x8m81_1/S pmos_1p2$$46284844_3v512x8m81
Xpmos_1p2$$46286892_3v512x8m81_0 vdd vdd nmos_5p04310591302028_3v512x8m81_1/S nmos_5p04310591302032_3v512x8m81_0/D
+ nmos_5p04310591302032_3v512x8m81_0/D nmos_5p04310591302032_3v512x8m81_0/D pmos_1p2$$46286892_3v512x8m81
Xnmos_5p04310591302023_3v512x8m81_0 vss pmos_5p04310591302027_3v512x8m81_2/S pmos_5p04310591302027_3v512x8m81_0/S
+ pmos_5p04310591302027_3v512x8m81_0/S vss nmos_5p04310591302023_3v512x8m81
Xnmos_5p04310591302028_3v512x8m81_1 nmos_5p04310591302028_3v512x8m81_1/D pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D nmos_5p04310591302028_3v512x8m81_1/S
+ pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D vss nmos_5p04310591302028_3v512x8m81
Xnmos_5p04310591302028_3v512x8m81_0 nmos_5p04310591302028_3v512x8m81_1/D nmos_5p04310591302032_3v512x8m81_0/D
+ nmos_5p04310591302032_3v512x8m81_0/D nmos_5p04310591302032_3v512x8m81_0/D nmos_5p04310591302032_3v512x8m81_0/D
+ vss nmos_5p04310591302032_3v512x8m81_0/D vss nmos_5p04310591302028_3v512x8m81
Xpmos_1p2$$46281772_3v512x8m81_0 vdd pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S
+ vdd pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81
Xpmos_1p2$$46281772_3v512x8m81_1 vdd pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S
+ nmos_5p04310591302028_3v512x8m81_1/S pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ vdd pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D pmos_1p2$$46281772_3v512x8m81
Xnmos_5p04310591302023_3v512x8m81_1 vss pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ vss pmos_5p04310591302027_3v512x8m81_1/S vss nmos_5p04310591302023_3v512x8m81
Xnmos_5p04310591302023_3v512x8m81_2 vss pmos_5p04310591302027_3v512x8m81_1/S pmos_5p04310591302027_3v512x8m81_2/S
+ pmos_5p04310591302027_3v512x8m81_2/S vss nmos_5p04310591302023_3v512x8m81
Xpmos_1p2$$46285868_3v512x8m81_0 vdd nmos_5p04310591302028_3v512x8m81_1/S pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ vdd pmos_1p2$$46285868_3v512x8m81
Xpmos_5p04310591302038_3v512x8m81_0 vdd pmos_5p04310591302027_3v512x8m81_0/S vdd pmos_5p04310591302038_3v512x8m81_0/S
+ pmos_5p04310591302038_3v512x8m81
Xnmos_1p2$$45103148_3v512x8m81_0 nmos_5p04310591302028_3v512x8m81_1/S pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D nmos_5p04310591302028_3v512x8m81_1/S
+ vss pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S vss nmos_1p2$$45103148_3v512x8m81
Xnmos_5p04310591302012_3v512x8m81_0 nmos_5p04310591302028_3v512x8m81_1/S se nmos_5p04310591302028_3v512x8m81_1/S
+ vss nmos_5p04310591302028_3v512x8m81_1/S nmos_5p04310591302028_3v512x8m81_1/S vss
+ nmos_5p04310591302012_3v512x8m81
Xpmos_1p2$$45095980_3v512x8m81_0 nmos_5p04310591302028_3v512x8m81_1/S nmos_5p04310591302028_3v512x8m81_1/S
+ nmos_5p04310591302028_3v512x8m81_1/S nmos_5p04310591302028_3v512x8m81_1/S se nmos_5p04310591302028_3v512x8m81_1/S
+ nmos_5p04310591302028_3v512x8m81_1/S nmos_5p04310591302028_3v512x8m81_1/S vdd nmos_5p04310591302028_3v512x8m81_1/S
+ nmos_5p04310591302028_3v512x8m81_1/S vdd nmos_5p04310591302028_3v512x8m81_1/S pmos_1p2$$45095980_3v512x8m81
Xpmos_5p04310591302027_3v512x8m81_0 vdd pmos_5p04310591302027_3v512x8m81_2/S pmos_5p04310591302027_3v512x8m81_0/S
+ vdd pmos_5p04310591302027_3v512x8m81_0/S pmos_5p04310591302027_3v512x8m81
Xpmos_1p2$$46282796_3v512x8m81_0 men vdd men men vdd pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ men men pmos_1p2$$46282796_3v512x8m81
Xpmos_5p04310591302027_3v512x8m81_1 vdd pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ vss vdd pmos_5p04310591302027_3v512x8m81_1/S pmos_5p04310591302027_3v512x8m81
Xnmos_1p2$$45100076_3v512x8m81_0 vss pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_1/pmos_5p04310591302025_3v512x8m81_0/S
+ vss nmos_1p2$$45100076_3v512x8m81
Xpmos_5p04310591302027_3v512x8m81_2 vdd pmos_5p04310591302027_3v512x8m81_1/S pmos_5p04310591302027_3v512x8m81_2/S
+ vdd pmos_5p04310591302027_3v512x8m81_2/S pmos_5p04310591302027_3v512x8m81
Xnmos_5p04310591302032_3v512x8m81_0 nmos_5p04310591302032_3v512x8m81_0/D pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D vss vss nmos_5p04310591302032_3v512x8m81
Xpmos_1p2$$46283820_3v512x8m81_0 pcb pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S vdd vdd pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S
+ pmos_1p2$$46281772_3v512x8m81_0/pmos_5p04310591302025_3v512x8m81_0/S pmos_1p2$$46283820_3v512x8m81
Xnmos_1p2$$45101100_3v512x8m81_0 men men vss men men pmos_1p2$$46282796_3v512x8m81_0/pmos_5p04310591302024_3v512x8m81_0/D
+ men vss nmos_1p2$$45101100_3v512x8m81
Xnmos_5p04310591302033_3v512x8m81_0 vss pmos_5p04310591302027_3v512x8m81_0/S pmos_5p04310591302038_3v512x8m81_0/S
+ vss nmos_5p04310591302033_3v512x8m81
Xpmos_1p2$$46287916_3v512x8m81_0 vdd pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D
+ vdd nmos_5p04310591302032_3v512x8m81_0/D pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D
+ pmos_1p2$$46287916_3v512x8m81
X0 pmos_1p2$$46284844_3v512x8m81_0/pmos_5p04310591302035_3v512x8m81_0/D pmos_5p04310591302027_3v512x8m81_1/S vss vss nfet_03v3 ad=0.2948p pd=2.22u as=0.2948p ps=2.22u w=0.67u l=0.28u
.ends

.subckt nmos_5p04310591302046_3v512x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X1 S a_662_n44# D VSUBS nfet_03v3 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.28u
X2 D a_502_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X3 S a_20_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X4 D a_181_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X5 D a_n140_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.28u
.ends

.subckt pmos_5p04310591302049_3v512x8m81 a_20_n44# D a_181_n44# a_n140_n44# S a_341_n44#
+ a_503_n44# a_663_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.4664p pd=2.29u as=0.4576p ps=2.28u w=1.76u l=0.28u
X1 S a_20_n44# D w_n314_n86# pfet_03v3 ad=0.462p pd=2.285u as=0.4576p ps=2.28u w=1.76u l=0.28u
X2 D a_181_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.462p ps=2.285u w=1.76u l=0.28u
X3 D a_n140_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.7744p ps=4.4u w=1.76u l=0.28u
X4 S a_663_n44# D w_n314_n86# pfet_03v3 ad=0.7832p pd=4.41u as=0.4576p ps=2.28u w=1.76u l=0.28u
X5 D a_503_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.4664p ps=2.29u w=1.76u l=0.28u
.ends

.subckt pmos_1p2$$171625516_3v512x8m81 a_n42_n34# pmos_5p0431059130203_3v512x8m81_0/w_n202_n86#
+ pmos_5p0431059130203_3v512x8m81_0/S a_118_n34# pmos_5p0431059130203_3v512x8m81_0/D
Xpmos_5p0431059130203_3v512x8m81_0 pmos_5p0431059130203_3v512x8m81_0/D a_n42_n34#
+ a_118_n34# pmos_5p0431059130203_3v512x8m81_0/w_n202_n86# pmos_5p0431059130203_3v512x8m81_0/S
+ pmos_5p0431059130203_3v512x8m81
.ends

.subckt nmos_5p04310591302050_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# VSUBS
X0 D a_265_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S a_104_n44# D VSUBS nfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302044_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.451p pd=2.93u as=0.451p ps=2.93u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302047_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.8206p pd=4.61u as=0.8206p ps=4.61u w=1.865u l=0.28u
.ends

.subckt nmos_5p04310591302045_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt pmos_5p04310591302048_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.924p pd=5.08u as=0.924p ps=5.08u w=2.1u l=0.28u
.ends

.subckt outbuf_oe_3v512x8m81 qp qn se q GWE vss vdd
Xpmos_5p04310591302013_3v512x8m81_0 pmos_5p04310591302013_3v512x8m81_0/D se pmos_5p04310591302051_3v512x8m81_0/D
+ se se vdd pmos_5p04310591302013_3v512x8m81
Xnmos_5p04310591302046_3v512x8m81_0 pmos_5p04310591302051_3v512x8m81_0/D vss pmos_5p04310591302051_3v512x8m81_0/D
+ pmos_5p04310591302051_3v512x8m81_0/D pmos_5p04310591302051_3v512x8m81_0/D pmos_5p04310591302051_3v512x8m81_0/D
+ q pmos_5p04310591302051_3v512x8m81_0/D vss nmos_5p04310591302046_3v512x8m81
Xpmos_5p04310591302049_3v512x8m81_0 pmos_5p04310591302051_3v512x8m81_0/D vdd pmos_5p04310591302051_3v512x8m81_0/D
+ pmos_5p04310591302051_3v512x8m81_0/D q pmos_5p04310591302051_3v512x8m81_0/D pmos_5p04310591302051_3v512x8m81_0/D
+ pmos_5p04310591302051_3v512x8m81_0/D vdd pmos_5p04310591302049_3v512x8m81
Xpmos_5p04310591302051_3v512x8m81_0 pmos_5p04310591302051_3v512x8m81_0/D qp qp vdd
+ pmos_5p04310591302051_3v512x8m81_1/S pmos_5p04310591302051_3v512x8m81
Xpmos_5p04310591302051_3v512x8m81_1 vdd pmos_5p04310591302048_3v512x8m81_0/S pmos_5p04310591302048_3v512x8m81_0/S
+ vdd pmos_5p04310591302051_3v512x8m81_1/S pmos_5p04310591302051_3v512x8m81
Xpmos_1p2$$171625516_3v512x8m81_0 pmos_5p04310591302038_3v512x8m81_0/D vdd vdd pmos_5p04310591302038_3v512x8m81_0/D
+ pmos_5p04310591302013_3v512x8m81_0/D pmos_1p2$$171625516_3v512x8m81
Xpmos_5p04310591302014_3v512x8m81_0 pmos_5p04310591302014_3v512x8m81_0/D se vdd vdd
+ pmos_5p04310591302014_3v512x8m81
Xpmos_5p04310591302038_3v512x8m81_0 pmos_5p04310591302038_3v512x8m81_0/D pmos_5p04310591302051_3v512x8m81_0/D
+ vdd vdd pmos_5p04310591302038_3v512x8m81
Xnmos_5p04310591302050_3v512x8m81_0 pmos_5p04310591302013_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_0/D
+ pmos_5p04310591302051_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_0/D pmos_5p04310591302014_3v512x8m81_0/D
+ vss nmos_5p04310591302050_3v512x8m81
Xnmos_5p04310591302044_3v512x8m81_0 vss pmos_5p04310591302047_3v512x8m81_0/S pmos_5p04310591302048_3v512x8m81_0/S
+ vss nmos_5p04310591302044_3v512x8m81
Xpmos_5p04310591302047_3v512x8m81_0 vdd GWE vdd pmos_5p04310591302047_3v512x8m81_0/S
+ pmos_5p04310591302047_3v512x8m81
Xnmos_5p04310591302033_3v512x8m81_0 pmos_5p04310591302038_3v512x8m81_0/D pmos_5p04310591302051_3v512x8m81_0/D
+ vss vss nmos_5p04310591302033_3v512x8m81
Xnmos_5p04310591302045_3v512x8m81_0 vss pmos_5p04310591302047_3v512x8m81_0/S pmos_5p04310591302047_3v512x8m81_0/S
+ nmos_5p04310591302045_3v512x8m81_1/S vss nmos_5p04310591302045_3v512x8m81
Xnmos_5p04310591302045_3v512x8m81_1 pmos_5p04310591302051_3v512x8m81_0/D qn qn nmos_5p04310591302045_3v512x8m81_1/S
+ vss nmos_5p04310591302045_3v512x8m81
Xpmos_5p04310591302048_3v512x8m81_0 vdd pmos_5p04310591302047_3v512x8m81_0/S vdd pmos_5p04310591302048_3v512x8m81_0/S
+ pmos_5p04310591302048_3v512x8m81
X0 vss pmos_5p04310591302038_3v512x8m81_0/D pmos_5p04310591302013_3v512x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss se pmos_5p04310591302014_3v512x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X2 pmos_5p04310591302047_3v512x8m81_0/S GWE vss vss nfet_03v3 ad=0.3278p pd=2.37u as=0.3278p ps=2.37u w=0.745u l=0.28u
.ends

.subckt saout_m2_3v512x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWEN GWE
+ bb[1] bb[3] bb[4] bb[5] bb[7] bb[6] b[5] b[6] b[7] b[2] q pcb b[1] b[3] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN din_3v512x8m81_0/men mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b bb[2] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb outbuf_oe_3v512x8m81_0/GWE mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass
+ ypass[7] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ b[4] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass vdd mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ vss mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
Xdin_3v512x8m81_0 vdd vdd vdd sa_3v512x8m81_0/wep din_3v512x8m81_0/men vdd vss vdd
+ pcb din_3v512x8m81
Xwen_wm1_3v512x8m81_0 GWEN din_3v512x8m81_0/men sa_3v512x8m81_0/wep WEN vdd vss wen_wm1_3v512x8m81
Xmux821_3v512x8m81_0 mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ vdd vdd vdd b[6] mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ bb[5] vdd vdd b[1] vdd mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ ypass[7] b[4] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb bb[3] vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ vdd vdd vss vdd pcb ypass[7] vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass b[3] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ bb[2] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass vss mux821_3v512x8m81
Xsa_3v512x8m81_0 sa_3v512x8m81_0/qp sa_3v512x8m81_0/wep sa_3v512x8m81_0/se pcb vdd
+ vss vdd sa_3v512x8m81
Xsacntl_2_3v512x8m81_0 pcb sa_3v512x8m81_0/se sacntl_2_3v512x8m81_0/pmos_5p04310591302027_3v512x8m81_2/S
+ sacntl_2_3v512x8m81_0/pmos_5p04310591302027_3v512x8m81_1/S din_3v512x8m81_0/men
+ vdd vss sacntl_2_3v512x8m81
Xoutbuf_oe_3v512x8m81_0 sa_3v512x8m81_0/qp sa_3v512x8m81_0/qp sa_3v512x8m81_0/se q
+ outbuf_oe_3v512x8m81_0/GWE vss vdd outbuf_oe_3v512x8m81
.ends

.subckt saout_R_m2_3v512x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWE GWEN
+ datain b[6] b[5] b[4] b[2] b[1] b[0] bb[6] bb[7] q bb[4] bb[3] bb[0] bb[1] pcb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b bb[2] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b WEN sa_3v512x8m81_0/pcb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ din_3v512x8m81_0/men mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ bb[5] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass ypass[7] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb m2_26_12231# mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ b[3] vdd vss mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
Xdin_3v512x8m81_0 vdd vdd datain sa_3v512x8m81_0/wep din_3v512x8m81_0/men vdd vss
+ vdd sa_3v512x8m81_0/pcb din_3v512x8m81
Xwen_wm1_3v512x8m81_0 GWEN din_3v512x8m81_0/men sa_3v512x8m81_0/wep WEN vdd vss wen_wm1_3v512x8m81
Xmux821_3v512x8m81_0 mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ vdd vdd vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ bb[2] vdd vdd b[6] vdd bb[7] vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/ypass b[3] ypass[7] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb bb[4] vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ vdd vdd m2_26_12231# vdd sa_3v512x8m81_0/pcb ypass[7] vdd mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/ypass vdd mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb bb[5] mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ vss mux821_3v512x8m81
Xsa_3v512x8m81_0 sa_3v512x8m81_0/qp sa_3v512x8m81_0/wep sa_3v512x8m81_0/se sa_3v512x8m81_0/pcb
+ vdd vss vdd sa_3v512x8m81
Xsacntl_2_3v512x8m81_0 sa_3v512x8m81_0/pcb sa_3v512x8m81_0/se sacntl_2_3v512x8m81_0/pmos_5p04310591302027_3v512x8m81_2/S
+ sacntl_2_3v512x8m81_0/pmos_5p04310591302027_3v512x8m81_1/S din_3v512x8m81_0/men
+ vdd vss sacntl_2_3v512x8m81
Xoutbuf_oe_3v512x8m81_0 sa_3v512x8m81_0/qp sa_3v512x8m81_0/qp sa_3v512x8m81_0/se q
+ GWE vss vdd outbuf_oe_3v512x8m81
.ends

.subckt col_512a_3v512x8m81 WL[3] ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] ypass[7]
+ WL[32] WL[30] WL[29] WL[22] WL[19] WL[49] WL[12] WL[11] WL[50] WL[51] WL[10] WL[43]
+ WL[35] WL[37] WL[7] WL[33] WL[6] WL[38] WL[36] WL[46] WL[55] WL[53] WL[17] WL[54]
+ WL[52] WL[16] WL[63] WL[14] WL[60] WL[13] WL[28] ypass[6] ypass[2] WL[25] b[1] b[7]
+ b[13] b[22] b[28] b[31] din[1] din[3] din[2] din[0] q[0] q[1] q[2] q[3] b[23] b[20]
+ b[14] b[11] b[8] bb[0] bb[1] bb[2] bb[9] bb[10] bb[11] bb[12] bb[13] bb[14] bb[15]
+ bb[19] bb[21] bb[22] bb[26] bb[28] bb[29] bb[31] b[30] b[27] b[12] b[0] b[3] b[18]
+ pcb[0] pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1] WEN[0] saout_R_m2_3v512x8m81_1/datain
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb WL[58] saout_m2_3v512x8m81_4/outbuf_oe_3v512x8m81_0/GWE
+ WL[0] saout_m2_3v512x8m81_4/GWEN saout_R_m2_3v512x8m81_0/datain saout_R_m2_3v512x8m81_0/q
+ m3_n771_22409# saout_m2_3v512x8m81_3/bb[2] WL[59] men WL[40] saout_m2_3v512x8m81_4/q
+ saout_R_m2_3v512x8m81_1/b[6] WL[23] saout_R_m2_3v512x8m81_0/GWE saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ WL[1] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[26] saout_m2_3v512x8m81_4/bb[5] WL[61] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[4] saout_m2_3v512x8m81_3/b[1] saout_m2_3v512x8m81_3/bb[3] saout_m2_3v512x8m81_3/b[4]
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb WL[56] saout_m2_3v512x8m81_4/GWE
+ saout_R_m2_3v512x8m81_1/b[3] WL[39] WL[20] WL[47] saout_m2_3v512x8m81_3/b[3] saout_R_m2_3v512x8m81_1/bb[7]
+ saout_m2_3v512x8m81_4/b[3] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_R_m2_3v512x8m81_0/bb[2]
+ bb[17] b[5] WL[41] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_m2_3v512x8m81_4/b[6] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[44] saout_m2_3v512x8m81_3/bb[5] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ WL[27] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb WL[5]
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb saout_R_m2_3v512x8m81_1/bb[4]
+ saout_R_m2_3v512x8m81_1/GWE WL[57] b[25] bb[8] WL[8] saout_R_m2_3v512x8m81_0/b[3]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ WL[21] saout_R_m2_3v512x8m81_1/bb[5] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b bb[6] WL[24]
+ GWE saout_R_m2_3v512x8m81_1/q WL[2] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_3/q b[10] WL[62] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb saout_m2_3v512x8m81_3/b[6]
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb WL[45] bb[24]
+ bb[4] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b WL[15] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[48] b[16] b[9] WL[18] saout_R_m2_3v512x8m81_0/bb[4] b[29] WL[31] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[9] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b WL[34]
+ bb[30] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb WL[42]
+ VDD saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b VSS
XCell_array8x8_3v512x8m81_0 saout_R_m2_3v512x8m81_1/b[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ saout_R_m2_3v512x8m81_1/b[3] b[5] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ saout_R_m2_3v512x8m81_1/bb[7] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ WL[58] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_m2_3v512x8m81_3/bb[2]
+ WL[29] bb[8] saout_R_m2_3v512x8m81_0/b[3] saout_R_m2_3v512x8m81_1/bb[4] WL[59] bb[6]
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_3/b[4] b[10] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb WL[35] saout_m2_3v512x8m81_3/b[3]
+ b[9] saout_R_m2_3v512x8m81_0/bb[4] WL[44] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ b[16] WL[20] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_m2_3v512x8m81_3/bb[5] WL[24] bb[11] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb WL[40] WL[50]
+ WL[49] saout_m2_3v512x8m81_4/bb[5] WL[54] b[25] WL[21] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb bb[10] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ bb[30] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b WL[51]
+ WL[48] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb saout_m2_3v512x8m81_3/b[1]
+ WL[45] WL[7] bb[17] bb[4] WL[31] WL[61] WL[17] WL[26] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ saout_m2_3v512x8m81_3/b[6] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ b[12] WL[47] bb[24] saout_R_m2_3v512x8m81_1/bb[5] WL[57] WL[0] WL[36] WL[46] WL[15]
+ WL[3] WL[56] saout_m2_3v512x8m81_4/b[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[25] saout_m2_3v512x8m81_3/bb[3] WL[14] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[22] WL[41] WL[2] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ b[29] WL[27] WL[4] WL[9] WL[12] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[18] WL[5] b[18] WL[52] WL[33] WL[13] WL[34] WL[55] saout_m2_3v512x8m81_4/b[3]
+ WL[32] VDD WL[30] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ WL[43] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb WL[28]
+ WL[63] WL[10] b[31] saout_R_m2_3v512x8m81_0/bb[2] WL[53] WL[6] WL[38] WL[62] WL[16]
+ WL[1] WL[39] WL[60] WL[37] WL[42] WL[8] WL[23] WL[19] WL[11] VSS Cell_array8x8_3v512x8m81
Xsaout_m2_3v512x8m81_4 saout_m2_3v512x8m81_4/ypass[2] saout_m2_3v512x8m81_4/ypass[3]
+ saout_m2_3v512x8m81_4/ypass[4] saout_m2_3v512x8m81_4/ypass[5] saout_m2_3v512x8m81_4/ypass[6]
+ saout_m2_3v512x8m81_4/GWEN saout_m2_3v512x8m81_4/GWE saout_m2_3v512x8m81_4/bb[1]
+ bb[11] saout_m2_3v512x8m81_4/bb[4] saout_m2_3v512x8m81_4/bb[5] saout_m2_3v512x8m81_4/bb[7]
+ saout_m2_3v512x8m81_4/bb[6] saout_m2_3v512x8m81_4/b[5] saout_m2_3v512x8m81_4/b[6]
+ saout_m2_3v512x8m81_4/b[7] saout_m2_3v512x8m81_4/b[2] saout_m2_3v512x8m81_4/q saout_m2_3v512x8m81_4/pcb
+ b[9] saout_m2_3v512x8m81_4/b[3] b[10] WEN[1] men saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b bb[10] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb saout_m2_3v512x8m81_4/outbuf_oe_3v512x8m81_0/GWE
+ ypass[6] ypass[5] ypass[7] ypass[2] ypass[0] saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb ypass[1] b[12]
+ ypass[4] VDD bb[8] VSS ypass[3] saout_m2_3v512x8m81
Xsaout_m2_3v512x8m81_3 saout_m2_3v512x8m81_3/ypass[2] saout_m2_3v512x8m81_3/ypass[3]
+ saout_m2_3v512x8m81_3/ypass[4] saout_m2_3v512x8m81_3/ypass[5] saout_m2_3v512x8m81_3/ypass[6]
+ saout_m2_3v512x8m81_4/GWEN GWE saout_m2_3v512x8m81_3/bb[1] saout_m2_3v512x8m81_3/bb[3]
+ saout_m2_3v512x8m81_3/bb[4] saout_m2_3v512x8m81_3/bb[5] saout_m2_3v512x8m81_3/bb[7]
+ saout_m2_3v512x8m81_3/bb[6] saout_m2_3v512x8m81_3/b[5] saout_m2_3v512x8m81_3/b[6]
+ saout_m2_3v512x8m81_3/b[7] saout_m2_3v512x8m81_3/b[2] saout_m2_3v512x8m81_3/q saout_m2_3v512x8m81_3/pcb
+ saout_m2_3v512x8m81_3/b[1] saout_m2_3v512x8m81_3/b[3] b[25] WEN[3] men saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ b[31] saout_m2_3v512x8m81_3/bb[2] b[29] bb[24] GWE ypass[6] ypass[5] ypass[7] ypass[2]
+ ypass[0] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb bb[30]
+ ypass[1] saout_m2_3v512x8m81_3/b[4] ypass[4] VDD saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ VSS ypass[3] saout_m2_3v512x8m81
Xsaout_R_m2_3v512x8m81_0 saout_R_m2_3v512x8m81_0/ypass[2] saout_R_m2_3v512x8m81_0/ypass[3]
+ saout_R_m2_3v512x8m81_0/ypass[4] saout_R_m2_3v512x8m81_0/ypass[5] saout_R_m2_3v512x8m81_0/ypass[6]
+ saout_R_m2_3v512x8m81_0/GWE saout_m2_3v512x8m81_4/GWEN saout_R_m2_3v512x8m81_0/datain
+ b[5] saout_R_m2_3v512x8m81_0/b[5] saout_R_m2_3v512x8m81_0/b[4] saout_R_m2_3v512x8m81_0/b[2]
+ saout_R_m2_3v512x8m81_0/b[1] saout_R_m2_3v512x8m81_0/b[0] saout_R_m2_3v512x8m81_0/bb[6]
+ bb[6] saout_R_m2_3v512x8m81_0/q saout_R_m2_3v512x8m81_0/bb[4] saout_R_m2_3v512x8m81_0/bb[3]
+ saout_R_m2_3v512x8m81_0/bb[0] saout_R_m2_3v512x8m81_0/bb[1] saout_R_m2_3v512x8m81_0/pcb
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_R_m2_3v512x8m81_0/bb[2] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b WEN[0] saout_R_m2_3v512x8m81_0/sa_3v512x8m81_0/pcb
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb men ypass[7]
+ ypass[6] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ bb[4] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb ypass[4]
+ saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b ypass[1] ypass[0]
+ ypass[5] ypass[2] saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ VSS saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb saout_R_m2_3v512x8m81_0/b[3]
+ VDD VSS ypass[3] saout_R_m2_3v512x8m81
Xsaout_R_m2_3v512x8m81_1 saout_R_m2_3v512x8m81_1/ypass[2] saout_R_m2_3v512x8m81_1/ypass[3]
+ saout_R_m2_3v512x8m81_1/ypass[4] saout_R_m2_3v512x8m81_1/ypass[5] saout_R_m2_3v512x8m81_1/ypass[6]
+ saout_R_m2_3v512x8m81_1/GWE saout_m2_3v512x8m81_4/GWEN saout_R_m2_3v512x8m81_1/datain
+ saout_R_m2_3v512x8m81_1/b[6] saout_R_m2_3v512x8m81_1/b[5] saout_R_m2_3v512x8m81_1/b[4]
+ saout_R_m2_3v512x8m81_1/b[2] saout_R_m2_3v512x8m81_1/b[1] saout_R_m2_3v512x8m81_1/b[0]
+ saout_R_m2_3v512x8m81_1/bb[6] saout_R_m2_3v512x8m81_1/bb[7] saout_R_m2_3v512x8m81_1/q
+ saout_R_m2_3v512x8m81_1/bb[4] saout_R_m2_3v512x8m81_1/bb[3] saout_R_m2_3v512x8m81_1/bb[0]
+ saout_R_m2_3v512x8m81_1/bb[1] saout_R_m2_3v512x8m81_1/pcb bb[17] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ b[18] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN[2] saout_R_m2_3v512x8m81_1/sa_3v512x8m81_0/pcb saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ men ypass[7] ypass[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_1/bb[5] b[16] ypass[4] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ ypass[1] ypass[0] ypass[5] ypass[2] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ VSS saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb saout_R_m2_3v512x8m81_1/b[3]
+ VDD VSS ypass[3] saout_R_m2_3v512x8m81
.ends

.subckt lcol4_512_3v512x8m81 WL[32] WL[33] WL[34] WL[38] WL[39] WL[35] WL[36] WL[37]
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[50] WL[51] WL[52] WL[53]
+ WL[54] WL[55] WL[56] WL[58] WL[60] WL[61] WL[62] WL[63] WL[25] WL[24] WL[23] WL[22]
+ WL[21] WL[20] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[8]
+ WL[6] WL[31] WL[30] WL[28] WL[27] WL[26] din[1] din[3] din[2] q[1] q[2] q[3] pcb[2]
+ pcb[3] pcb[0] pcb[1] WEN[3] WEN[2] WEN[1] WEN[0] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/q
+ col_512a_3v512x8m81_0/WL[40] col_512a_3v512x8m81_0/WL[41] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/datain
+ col_512a_3v512x8m81_0/WL[43] col_512a_3v512x8m81_0/WL[60] WL[59] col_512a_3v512x8m81_0/WL[45]
+ col_512a_3v512x8m81_0/WL[62] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/GWE col_512a_3v512x8m81_0/WL[47]
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/outbuf_oe_3v512x8m81_0/GWE col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/GWEN
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/GWE col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/q
+ WL[0] col_512a_3v512x8m81_0/WL[10] col_512a_3v512x8m81_0/men WL[1] WL[2] col_512a_3v512x8m81_0/WL[12]
+ WL[3] col_512a_3v512x8m81_0/WL[13] WL[29] WL[4] col_512a_3v512x8m81_0/WL[14] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/q
+ WL[5] col_512a_3v512x8m81_0/WL[15] col_512a_3v512x8m81_0/WL[32] col_512a_3v512x8m81_0/WL[6]
+ WL[48] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/GWE WL[7] col_512a_3v512x8m81_0/WL[17]
+ col_512a_3v512x8m81_0/WL[34] col_512a_3v512x8m81_0/ypass[0] WL[49] col_512a_3v512x8m81_0/WL[8]
+ col_512a_3v512x8m81_0/ypass[1] WL[9] col_512a_3v512x8m81_0/WL[19] col_512a_3v512x8m81_0/WL[36]
+ col_512a_3v512x8m81_0/ypass[2] col_512a_3v512x8m81_0/ypass[3] col_512a_3v512x8m81_0/WL[38]
+ col_512a_3v512x8m81_0/ypass[4] col_512a_3v512x8m81_0/WL[39] col_512a_3v512x8m81_0/ypass[5]
+ col_512a_3v512x8m81_0/ypass[6] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/q col_512a_3v512x8m81_0/ypass[7]
+ col_512a_3v512x8m81_0/WL[58] WL[57] col_512a_3v512x8m81_0/GWE col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/datain
+ WL[19] VDD VSUBS col_512a_3v512x8m81_0/WL[21]
Xldummy_3v512x4_3v512x8m81_0 VSUBS VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[6] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[2]
+ col_512a_3v512x8m81_0/WL[32] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/bb[5] VDD
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[4] col_512a_3v512x8m81_0/b[25]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[3] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[3]
+ WL[32] VDD col_512a_3v512x8m81_0/WL[14] VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[6] WL[53] VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[3]
+ VDD WL[50] VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[3] col_512a_3v512x8m81_0/WL[17]
+ VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[4] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ VDD col_512a_3v512x8m81_0/b[12] col_512a_3v512x8m81_0/WL[34] VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ col_512a_3v512x8m81_0/bb[4] col_512a_3v512x8m81_0/b[29] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[5]
+ col_512a_3v512x8m81_0/WL[12] WL[36] VDD VSUBS VSUBS VDD VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/bb[6] WL[55] VSUBS VDD col_512a_3v512x8m81_0/b[29] WL[48]
+ VDD VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[5] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[5] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ VDD WL[29] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[6] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/b[3]
+ VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[6] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[4] col_512a_3v512x8m81_0/WL[10] col_512a_3v512x8m81_0/WL[39]
+ VSUBS VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/b[5] VDD WL[57] VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ VDD WL[46] VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[4] WL[30] VSUBS
+ VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[4] VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[27] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[2] VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ col_512a_3v512x8m81_0/WL[8] VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[4]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ col_512a_3v512x8m81_0/bb[30] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[6] WL[61]
+ VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ col_512a_3v512x8m81_0/bb[6] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[5] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[3] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/WL[19] VSUBS VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ col_512a_3v512x8m81_0/bb[30] col_512a_3v512x8m81_0/bb[4] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[6]
+ col_512a_3v512x8m81_0/WL[41] VSUBS VDD WL[59] VDD col_512a_3v512x8m81_0/b[31] VSUBS
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[1] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[3] VDD WL[44] VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/b[18] VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ WL[25] VDD col_512a_3v512x8m81_0/WL[21] VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/b[3]
+ VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ VDD col_512a_3v512x8m81_0/WL[43] col_512a_3v512x8m81_0/WL[6] VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ VDD WL[3] VSUBS VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[7] WL[5] VSUBS
+ col_512a_3v512x8m81_0/bb[8] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/b[18] WL[42] VDD VSUBS col_512a_3v512x8m81_0/bb[8] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/bb[17] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[22] VDD WL[23] VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[2]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ WL[4] col_512a_3v512x8m81_0/WL[45] VSUBS VSUBS col_512a_3v512x8m81_0/WL[62] VDD
+ VSUBS WL[7] VSUBS col_512a_3v512x8m81_0/b[9] VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/bb[17] VDD WL[40] VSUBS col_512a_3v512x8m81_0/b[9] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/b[16] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[21] WL[24] VDD VSUBS VSUBS VDD col_512a_3v512x8m81_0/WL[47] WL[0] VSUBS VSUBS
+ VDD col_512a_3v512x8m81_0/WL[60] VSUBS VDD WL[9] VSUBS col_512a_3v512x8m81_0/bb[10]
+ col_512a_3v512x8m81_0/b[10] col_512a_3v512x8m81_0/b[16] VDD col_512a_3v512x8m81_0/WL[40]
+ VDD VSUBS col_512a_3v512x8m81_0/bb[10] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/b[10] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[26] WL[19] VSUBS VDD VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[3]
+ col_512a_3v512x8m81_0/bb[11] WL[2] WL[47] VSUBS VSUBS col_512a_3v512x8m81_0/WL[58]
+ VDD VSUBS WL[11] col_512a_3v512x8m81_0/b[31] VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ VDD col_512a_3v512x8m81_0/WL[38] VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[1] col_512a_3v512x8m81_0/bb[24] WL[17]
+ WL[28] VDD VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/bb[5] WL[49] VSUBS VDD WL[54] VDD VSUBS
+ col_512a_3v512x8m81_0/WL[13] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[3] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[7]
+ VDD col_512a_3v512x8m81_0/WL[36] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[1]
+ col_512a_3v512x8m81_0/bb[11] VDD VSUBS col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/bb[24] col_512a_3v512x8m81_0/b[5] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[2]
+ col_512a_3v512x8m81_0/b[25] VDD WL[15] WL[34] VDD VSUBS VSUBS VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/b[12] WL[51] VSUBS VDD VDD VSUBS WL[52] VDD VSUBS VDD col_512a_3v512x8m81_0/WL[15]
+ ldummy_3v512x4_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[0] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[1] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[2] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[3] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[4] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[5] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[6] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[7] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[8] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[9] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[10] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[11] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[12] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[13] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[14] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[15] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[16] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[17] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[18] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[19] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[20] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[21] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[22] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[23] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[24] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[25] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[26] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[27] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[28] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[29] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[30] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[31] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[32] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[33] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[34] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[35] VDD VSUBS VDD dcap_103_novia_3v512x8m81
Xcol_512a_3v512x8m81_0 WL[3] col_512a_3v512x8m81_0/ypass[0] col_512a_3v512x8m81_0/ypass[1]
+ col_512a_3v512x8m81_0/ypass[3] col_512a_3v512x8m81_0/ypass[4] col_512a_3v512x8m81_0/ypass[5]
+ col_512a_3v512x8m81_0/ypass[7] col_512a_3v512x8m81_0/WL[32] WL[29] WL[28] WL[21]
+ col_512a_3v512x8m81_0/WL[19] WL[47] col_512a_3v512x8m81_0/WL[12] WL[11] WL[48] WL[49]
+ col_512a_3v512x8m81_0/WL[10] col_512a_3v512x8m81_0/WL[43] WL[34] WL[36] WL[7] WL[32]
+ col_512a_3v512x8m81_0/WL[6] col_512a_3v512x8m81_0/WL[38] col_512a_3v512x8m81_0/WL[36]
+ WL[44] WL[53] WL[51] col_512a_3v512x8m81_0/WL[17] WL[52] WL[50] WL[15] WL[61] col_512a_3v512x8m81_0/WL[14]
+ col_512a_3v512x8m81_0/WL[60] col_512a_3v512x8m81_0/WL[13] WL[27] col_512a_3v512x8m81_0/ypass[6]
+ col_512a_3v512x8m81_0/ypass[2] WL[24] col_512a_3v512x8m81_0/b[1] col_512a_3v512x8m81_0/b[7]
+ col_512a_3v512x8m81_0/b[13] col_512a_3v512x8m81_0/b[22] col_512a_3v512x8m81_0/b[28]
+ col_512a_3v512x8m81_0/b[31] col_512a_3v512x8m81_0/din[1] col_512a_3v512x8m81_0/din[3]
+ col_512a_3v512x8m81_0/din[2] col_512a_3v512x8m81_0/din[0] col_512a_3v512x8m81_0/q[0]
+ col_512a_3v512x8m81_0/q[1] col_512a_3v512x8m81_0/q[2] col_512a_3v512x8m81_0/q[3]
+ col_512a_3v512x8m81_0/b[23] col_512a_3v512x8m81_0/b[20] col_512a_3v512x8m81_0/b[14]
+ col_512a_3v512x8m81_0/b[11] col_512a_3v512x8m81_0/b[8] col_512a_3v512x8m81_0/bb[0]
+ col_512a_3v512x8m81_0/bb[1] col_512a_3v512x8m81_0/bb[2] col_512a_3v512x8m81_0/bb[9]
+ col_512a_3v512x8m81_0/bb[10] col_512a_3v512x8m81_0/bb[11] col_512a_3v512x8m81_0/bb[12]
+ col_512a_3v512x8m81_0/bb[13] col_512a_3v512x8m81_0/bb[14] col_512a_3v512x8m81_0/bb[15]
+ col_512a_3v512x8m81_0/bb[19] col_512a_3v512x8m81_0/bb[21] col_512a_3v512x8m81_0/bb[22]
+ col_512a_3v512x8m81_0/bb[26] col_512a_3v512x8m81_0/bb[28] col_512a_3v512x8m81_0/bb[29]
+ col_512a_3v512x8m81_0/bb[31] col_512a_3v512x8m81_0/b[30] col_512a_3v512x8m81_0/b[27]
+ col_512a_3v512x8m81_0/b[12] col_512a_3v512x8m81_0/b[0] col_512a_3v512x8m81_0/b[3]
+ col_512a_3v512x8m81_0/b[18] col_512a_3v512x8m81_0/pcb[0] col_512a_3v512x8m81_0/pcb[1]
+ col_512a_3v512x8m81_0/pcb[3] col_512a_3v512x8m81_0/pcb[2] WEN[3] WEN[2] WEN[1] WEN[0]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/datain col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/WL[58] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/outbuf_oe_3v512x8m81_0/GWE
+ WL[0] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/GWEN col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/datain
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/q VSUBS col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[2]
+ WL[57] col_512a_3v512x8m81_0/men col_512a_3v512x8m81_0/WL[40] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/q
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[6] WL[22] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/GWE
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ WL[1] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[25] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/bb[5] WL[59] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[4] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[1] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[3]
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[4] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[54] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/GWE col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/b[3]
+ col_512a_3v512x8m81_0/WL[39] WL[19] col_512a_3v512x8m81_0/WL[47] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[3]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[7] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[3]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[2] col_512a_3v512x8m81_0/bb[17]
+ col_512a_3v512x8m81_0/b[5] col_512a_3v512x8m81_0/WL[41] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/b[6] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[42] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/bb[5] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ WL[26] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[5] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[4] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/GWE
+ WL[55] col_512a_3v512x8m81_0/b[25] col_512a_3v512x8m81_0/bb[8] col_512a_3v512x8m81_0/WL[8]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/b[3] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/WL[21] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/bb[5]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ col_512a_3v512x8m81_0/bb[6] WL[23] col_512a_3v512x8m81_0/GWE col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/q
+ WL[2] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/q col_512a_3v512x8m81_0/b[10] col_512a_3v512x8m81_0/WL[62]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/b[6] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ col_512a_3v512x8m81_0/WL[45] col_512a_3v512x8m81_0/bb[24] col_512a_3v512x8m81_0/bb[4]
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ col_512a_3v512x8m81_0/WL[15] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[46] col_512a_3v512x8m81_0/b[16] col_512a_3v512x8m81_0/b[9] WL[17] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/bb[4]
+ col_512a_3v512x8m81_0/b[29] WL[30] col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ col_512a_3v512x8m81_0/saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[9] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ col_512a_3v512x8m81_0/WL[34] col_512a_3v512x8m81_0/bb[30] col_512a_3v512x8m81_0/saout_R_m2_3v512x8m81_0/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[40] VDD col_512a_3v512x8m81_0/saout_m2_3v512x8m81_4/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ VSUBS col_512a_3v512x8m81
.ends

.subckt nmos_5p04310591302096_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=1.0309p pd=4.485u as=1.7446p ps=8.81u w=3.965u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=1.7446p pd=8.81u as=1.0309p ps=4.485u w=3.965u l=0.28u
.ends

.subckt x018SRAM_cell1_dummy_R_3v512x8m81 m3_82_330# a_248_342# a_62_178# w_30_512#
+ a_430_96# a_110_96# a_192_298# VSUBS
X0 a_192_298# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_408_342# a_248_342# a_192_298# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_408_342# a_248_342# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_408_342# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt ypass_gate_3v512x8m81_0 bb db ypass d pcb m3_0_2091# m3_0_2831# pmos_5p0431059130201_3v512x8m81_2/D
+ a_64_1295# m3_0_3056# pmos_5p0431059130201_3v512x8m81_0/D m3_0_3781# vdd m3_0_1632#
+ vss m3_0_3536# m3_0_3291# b m3_0_2331# m3_0_2581#
Xnmos_5p0431059130200_3v512x8m81_0 pmos_5p0431059130201_3v512x8m81_2/D a_64_1295#
+ bb vss nmos_5p0431059130200_3v512x8m81
Xnmos_5p0431059130200_3v512x8m81_1 pmos_5p0431059130201_3v512x8m81_0/D a_64_1295#
+ b vss nmos_5p0431059130200_3v512x8m81
Xnmos_5p0431059130202_3v512x8m81_0 nmos_5p0431059130202_3v512x8m81_0/D a_64_1295#
+ a_64_1295# vss vss nmos_5p0431059130202_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_0 pmos_5p0431059130201_3v512x8m81_0/D nmos_5p0431059130202_3v512x8m81_0/D
+ vdd b pmos_5p0431059130201_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_1 b pcb vdd bb pmos_5p0431059130201_3v512x8m81
Xpmos_5p0431059130201_3v512x8m81_2 pmos_5p0431059130201_3v512x8m81_2/D nmos_5p0431059130202_3v512x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v512x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
X1 bb pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X2 nmos_5p0431059130202_3v512x8m81_0/D a_64_1295# vdd vdd pfet_03v3 ad=0.1946p pd=1.255u as=0.38225p ps=2.49u w=0.695u l=0.28u
X3 vdd a_64_1295# nmos_5p0431059130202_3v512x8m81_0/D vdd pfet_03v3 ad=0.50735p pd=2.85u as=0.1946p ps=1.255u w=0.695u l=0.28u
X4 b pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X5 vdd pcb bb vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
.ends

.subckt pmos_5p04310591302095_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4251p pd=2.155u as=0.7194p ps=4.15u w=1.635u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7194p pd=4.15u as=0.4251p ps=2.155u w=1.635u l=0.28u
.ends

.subckt nmos_5p04310591302098_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1664p pd=1.16u as=0.2816p ps=2.16u w=0.64u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.2816p pd=2.16u as=0.1664p ps=1.16u w=0.64u l=0.28u
.ends

.subckt pmos_5p04310591302097_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.2909p pd=5.485u as=2.1846p ps=10.81u w=4.965u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=2.1846p pd=10.81u as=1.2909p ps=5.485u w=4.965u l=0.28u
.ends

.subckt rdummy_3v512x4_3v512x8m81 018SRAM_cell1_dummy_3v512x8m81_56/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_17/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_56/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_17/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_42/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_8/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_42/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_27/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/a_248_342# pmos_5p04310591302097_3v512x8m81_0/D
+ 018SRAM_cell1_dummy_3v512x8m81_27/m2_134_89# m3_15667_n5798# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_13/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_13/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_2/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_2/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_7/a_192_298# 018SRAM_cell1_dummy_R_3v512x8m81_55/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_64/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_37/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_37/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_62/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_23/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_62/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_23/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_65/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_47/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_47/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_33/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/a_248_342# w_15880_n13729#
+ 018SRAM_cell1_dummy_R_3v512x8m81_33/a_248_342# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v512x8m81_36/a_192_298# 018SRAM_cell1_dummy_3v512x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_57/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_57/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_18/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_43/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_43/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_55/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_28/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_28/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_53/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_14/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/w_30_512# ypass_gate_3v512x8m81_0_0/pcb
+ 018SRAM_cell1_dummy_R_3v512x8m81_53/a_248_342# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_3/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_14/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_56/a_192_298# 018SRAM_cell1_dummy_R_3v512x8m81_3/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_5/a_192_298# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_38/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_38/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_24/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_63/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_63/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_24/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_48/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_48/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_36/w_30_512# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ m1_16100_n16182# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_34/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_34/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_37/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_19/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_19/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_44/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_44/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_32/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_65/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_29/m2_346_89# ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D
+ 018SRAM_cell1_dummy_3v512x8m81_29/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_54/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_15/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_54/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_15/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_57/a_192_298#
+ 018SRAM_cell1_dummy_R_3v512x8m81_4/a_248_342# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v512x8m81_3/a_192_298# 018SRAM_cell1_dummy_R_3v512x8m81_61/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_39/m2_346_89# 018SRAM_cell1_dummy_R_3v512x8m81_5/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_39/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_64/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_25/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_64/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_25/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/m3_82_330# pmos_5p04310591302097_3v512x8m81_0/S
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_49/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_49/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_6/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_35/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_35/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_38/a_192_298# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_59/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_59/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_45/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_45/a_248_342# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_55/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_16/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_55/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_5/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_16/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_5/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_58/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_65/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_65/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_26/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_56/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_36/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_36/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_39/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# m3_15667_n5552# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_46/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_46/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_20/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_20/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_56/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_17/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_56/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_17/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_6/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_30/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_37/w_30_512# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_30/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_27/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_27/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_40/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_40/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_33/w_30_512# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_37/m3_82_330# m3_15667_n6510# 018SRAM_cell1_dummy_R_3v512x8m81_37/a_248_342#
+ pmos_5p04310591302095_3v512x8m81_0/S 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_50/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_50/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_47/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_62/w_30_512# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_47/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_3/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_60/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_60/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_21/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_18/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_57/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_57/a_248_342# 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_7/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_18/a_248_342#
+ m3_15667_n6288# 018SRAM_cell1_dummy_R_3v512x8m81_7/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_0/a_192_298#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89# 018SRAM_cell1_dummy_R_3v512x8m81_2/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89#
+ ypass_gate_3v512x8m81_0_0/vdd 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v512x8m81_28/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_28/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_41/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/a_248_342# a_16524_38786#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_41/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_38/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_38/a_248_342# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_51/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_48/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_48/a_248_342# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_40/a_192_298# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v512x8m81_61/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_22/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_0/a_248_342# m3_15698_n15942#
+ 018SRAM_cell1_dummy_3v512x8m81_61/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_22/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_58/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_58/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_8/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_8/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_1/a_192_298#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_32/m2_346_89# 018SRAM_cell1_dummy_R_3v512x8m81_57/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# m3_15667_n7247# 018SRAM_cell1_dummy_3v512x8m81_32/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_29/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_29/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_60/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_42/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_53/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_42/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_39/a_248_342# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_31/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_52/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_52/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_49/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_49/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_38/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_64/a_192_298# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_62/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_23/m2_346_89#
+ a_16524_2# 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_62/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_23/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_59/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_59/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_9/a_248_342# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v512x8m81_8/a_192_298# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_33/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_34/w_30_512# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_33/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_61/a_192_298#
+ 018SRAM_cell1_dummy_3v512x8m81_43/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_43/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_63/w_30_512#
+ m3_15645_n13711# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_32/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_53/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_53/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_4/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_63/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_24/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_63/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_24/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_10/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_10/a_248_342# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_6/a_192_298# 018SRAM_cell1_dummy_R_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_34/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v512x8m81_34/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_20/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_20/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_62/a_192_298# ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_3v512x8m81_44/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_40/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_44/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_30/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_30/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_33/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_54/m2_346_89# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_dummy_3v512x8m81_54/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_40/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_40/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_58/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_64/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_25/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_25/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_64/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_50/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_50/a_248_342# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_11/a_248_342# m3_15667_n6043# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_53/a_192_298#
+ 018SRAM_cell1_dummy_R_3v512x8m81_2/a_192_298# 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_35/m2_346_89# 018SRAM_cell1_dummy_R_3v512x8m81_54/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_35/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_60/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v512x8m81_21/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_60/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_21/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_63/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_dummy_3v512x8m81_45/m2_346_89#
+ 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v512x8m81_45/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v512x8m81_31/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_39/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v512x8m81_31/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_34/a_192_298#
+ 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_16/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_16/m2_134_89#
+ 018SRAM_cell1_dummy_3v512x8m81_55/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v512x8m81_41/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_41/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_35/w_30_512# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v512x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_26/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_51/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_12/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_51/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_12/a_248_342# 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_54/a_192_298# 018SRAM_cell1_dummy_R_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_4/a_192_298# 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89# 018SRAM_cell1_dummy_R_3v512x8m81_31/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_36/m2_346_89# 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89#
+ 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ m3_15667_n7002# 018SRAM_cell1_dummy_3v512x8m81_36/m2_134_89# 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_22/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_61/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_61/a_248_342# a_n547_48# 018SRAM_cell1_dummy_R_3v512x8m81_22/a_248_342#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v512x8m81_46/m2_346_89# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v512x8m81_60/w_30_512#
+ 018SRAM_cell1_dummy_3v512x8m81_46/m2_134_89# 018SRAM_cell1_dummy_R_3v512x8m81_7/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v512x8m81_32/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v512x8m81_32/a_248_342# 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v512x8m81_35/a_192_298#
+ m3_15667_n6752#
X018SRAM_cell1_dummy_3v512x8m81_6 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_6/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_7 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_7/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_8 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_8/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_9 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_9/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_30 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_0/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_20 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_20/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_31 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
Xnmos_5p04310591302096_3v512x8m81_0 pmos_5p04310591302097_3v512x8m81_0/D pmos_5p04310591302095_3v512x8m81_0/D
+ pmos_5p04310591302095_3v512x8m81_0/D ypass_gate_3v512x8m81_0_0/vss ypass_gate_3v512x8m81_0_0/vss
+ nmos_5p04310591302096_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_1/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_10 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_10/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_21 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_21/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_60 018SRAM_cell1_dummy_R_3v512x8m81_60/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_60/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_60/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_60/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_2/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_11 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_11/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_22 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_22/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_0 018SRAM_cell1_dummy_R_3v512x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_0/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_0/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_0/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_61 018SRAM_cell1_dummy_R_3v512x8m81_61/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_61/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_61/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_61/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_50 018SRAM_cell1_dummy_R_3v512x8m81_50/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_50/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_60/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_60/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_3/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_12 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_12/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_23 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96#
+ ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_1 018SRAM_cell1_dummy_R_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_1/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_1/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_1/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_62 018SRAM_cell1_dummy_R_3v512x8m81_62/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_62/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_62/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_62/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_51 018SRAM_cell1_dummy_R_3v512x8m81_51/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_51/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_58/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_58/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_40 018SRAM_cell1_dummy_R_3v512x8m81_40/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_40/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_40/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_40/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_4 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_4/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_13 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_13/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_24 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_24/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_2 018SRAM_cell1_dummy_R_3v512x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_2/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_2/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_2/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_63 018SRAM_cell1_dummy_R_3v512x8m81_63/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_63/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_63/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_63/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_52 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss
+ a_16524_38786# 018SRAM_cell1_3v512x8m81_1/w_30_512# ypass_gate_3v512x8m81_0_0/bb
+ ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_3v512x8m81_1/w_30_512# ypass_gate_3v512x8m81_0_0/vss
+ x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_41 018SRAM_cell1_dummy_R_3v512x8m81_41/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_41/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_64/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_64/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_30 018SRAM_cell1_dummy_R_3v512x8m81_30/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_30/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_39/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_39/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_5 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_5/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_3 018SRAM_cell1_dummy_R_3v512x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_3/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_3/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_3/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_14 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_31/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_14/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_25 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_30/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_25/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_60 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_60/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_60/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_64 018SRAM_cell1_dummy_R_3v512x8m81_64/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_64/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_64/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_64/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_53 018SRAM_cell1_dummy_R_3v512x8m81_53/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_53/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_53/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_53/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_42 018SRAM_cell1_dummy_R_3v512x8m81_42/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_42/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_53/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_53/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_31 018SRAM_cell1_dummy_R_3v512x8m81_31/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_31/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_31/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_31/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_20 018SRAM_cell1_dummy_R_3v512x8m81_20/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_20/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_31/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_31/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_6 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_15 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_15/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_26 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_26/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_50 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_50/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_61 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_61/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_61/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_4 018SRAM_cell1_dummy_R_3v512x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_4/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_4/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_4/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_65 018SRAM_cell1_dummy_R_3v512x8m81_65/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_65/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_65/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_65/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_54 018SRAM_cell1_dummy_R_3v512x8m81_54/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_54/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_54/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_54/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_43 018SRAM_cell1_dummy_R_3v512x8m81_43/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_43/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_57/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_57/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_32 018SRAM_cell1_dummy_R_3v512x8m81_32/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_32/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_32/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_32/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_21 018SRAM_cell1_dummy_R_3v512x8m81_21/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_21/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_35/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_35/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_10 018SRAM_cell1_dummy_R_3v512x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_10/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_0/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_0/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_7 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_7/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_5 018SRAM_cell1_dummy_R_3v512x8m81_5/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_5/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_5/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_5/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_16 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_16/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_27 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_27/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_40 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_40/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_40/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_51 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_51/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_62 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_62/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_62/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
Xypass_gate_3v512x8m81_0_0 ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/db
+ ypass_gate_3v512x8m81_0_0/ypass ypass_gate_3v512x8m81_0_0/d ypass_gate_3v512x8m81_0_0/pcb
+ m3_15667_n7247# m3_15667_n6510# ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/vdd
+ m3_15667_n6288# ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D m3_15667_n5552#
+ ypass_gate_3v512x8m81_0_0/vdd ypass_gate_3v512x8m81_0_0/vdd ypass_gate_3v512x8m81_0_0/vss
+ m3_15667_n5798# m3_15667_n6043# ypass_gate_3v512x8m81_0_0/b m3_15667_n7002# m3_15667_n6752#
+ ypass_gate_3v512x8m81_0
X018SRAM_cell1_dummy_R_3v512x8m81_55 018SRAM_cell1_dummy_R_3v512x8m81_55/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_55/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_55/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_55/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_44 018SRAM_cell1_dummy_R_3v512x8m81_44/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_44/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_55/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_55/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_33 018SRAM_cell1_dummy_R_3v512x8m81_33/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_33/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_33/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_33/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_22 018SRAM_cell1_dummy_R_3v512x8m81_22/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_22/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_37/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_37/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_11 018SRAM_cell1_dummy_R_3v512x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_11/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_1/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_1/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_8 a_n547_1214# 018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_0/m3_82_330# a_n547_1214#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96#
+ ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96# x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_17 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_17/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_28 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_28/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_30 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_30/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_41 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_41/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_41/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_52 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_52/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_52/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_63 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_63/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_63/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_6 018SRAM_cell1_dummy_R_3v512x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_6/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_6/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_6/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_56 018SRAM_cell1_dummy_R_3v512x8m81_56/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_56/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_56/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_56/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_45 018SRAM_cell1_dummy_R_3v512x8m81_45/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_45/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_62/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_62/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_34 018SRAM_cell1_dummy_R_3v512x8m81_34/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_34/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_34/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_34/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_23 018SRAM_cell1_dummy_R_3v512x8m81_23/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_23/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_36/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_36/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_12 018SRAM_cell1_dummy_R_3v512x8m81_12/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_12/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_8/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_8/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_9 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
Xpmos_5p04310591302095_3v512x8m81_0 pmos_5p04310591302095_3v512x8m81_0/D ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D pmos_5p04310591302095_3v512x8m81_0/S
+ pmos_5p04310591302095_3v512x8m81_0/S pmos_5p04310591302095_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_7 018SRAM_cell1_dummy_R_3v512x8m81_7/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_7/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_7/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_7/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_18 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_18/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/a_248_592# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_29 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_29/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_20 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_20/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_31 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_31/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_42 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_42/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_42/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_53 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_53/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_53/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_64 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_64/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_57 018SRAM_cell1_dummy_R_3v512x8m81_57/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_57/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_57/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_57/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_46 018SRAM_cell1_dummy_R_3v512x8m81_46/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_46/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_54/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_54/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_35 018SRAM_cell1_dummy_R_3v512x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_35/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_35/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_35/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_24 018SRAM_cell1_dummy_R_3v512x8m81_24/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_24/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_32/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_32/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_13 018SRAM_cell1_dummy_R_3v512x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_13/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_6/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_6/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_19 a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/a_248_342# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/m3_82_330#
+ a_n547_1214# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/a_248_342# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/a_248_592# 018SRAM_cell1_2x_3v512x8m81_19/018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/a_430_96# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_8 018SRAM_cell1_dummy_R_3v512x8m81_8/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_8/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_8/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_8/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_10 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_10/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_21 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_21/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_32 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_32/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_32/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_43 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_43/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_43/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_54 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_54/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_54/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_58 018SRAM_cell1_dummy_R_3v512x8m81_58/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_58/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_58/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_58/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_47 018SRAM_cell1_dummy_R_3v512x8m81_47/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_47/a_248_342# a_16524_38786# 018SRAM_cell1_dummy_R_3v512x8m81_56/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_56/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_36 018SRAM_cell1_dummy_R_3v512x8m81_36/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_36/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_36/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_36/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_25 018SRAM_cell1_dummy_R_3v512x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_25/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_33/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_33/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_14 018SRAM_cell1_dummy_R_3v512x8m81_14/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_14/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_2/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_2/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_11 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_11/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_22 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_22/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_33 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_33/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_33/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_44 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_44/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_44/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_55 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_55/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_9 018SRAM_cell1_dummy_R_3v512x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_9/a_248_342# a_16524_2# 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_59 018SRAM_cell1_dummy_R_3v512x8m81_59/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_59/a_248_342# a_16524_38786# 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_48 018SRAM_cell1_dummy_R_3v512x8m81_48/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_48/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_61/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_61/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_37 018SRAM_cell1_dummy_R_3v512x8m81_37/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_37/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_37/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_37/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_26 018SRAM_cell1_dummy_R_3v512x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_26/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_65/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_65/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_15 018SRAM_cell1_dummy_R_3v512x8m81_15/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_15/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_4/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_4/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_12 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_12/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_23 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_23/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_34 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_34/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_34/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_45 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_45/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_56 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_56/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_49 018SRAM_cell1_dummy_R_3v512x8m81_49/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_49/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_63/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_63/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_38 018SRAM_cell1_dummy_R_3v512x8m81_38/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_38/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_38/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_38/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_27 018SRAM_cell1_dummy_R_3v512x8m81_27/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_27/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_38/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_38/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_16 018SRAM_cell1_dummy_R_3v512x8m81_16/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_16/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_7/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_7/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_13 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_13/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_24 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_24/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_35 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_35/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_35/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_46 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_46/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_57 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_57/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_57/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_39 018SRAM_cell1_dummy_R_3v512x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_39/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_39/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_39/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_28 018SRAM_cell1_dummy_R_3v512x8m81_28/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_28/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_40/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_40/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_17 018SRAM_cell1_dummy_R_3v512x8m81_17/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_17/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_5/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_5/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_14 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_14/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_25 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_25/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_36 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_36/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_36/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_47 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_47/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_47/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_29 018SRAM_cell1_dummy_R_3v512x8m81_29/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_29/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_34/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_34/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_18 018SRAM_cell1_dummy_R_3v512x8m81_18/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v512x8m81_18/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v512x8m81_3/w_30_512#
+ ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b 018SRAM_cell1_dummy_R_3v512x8m81_3/a_192_298#
+ ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
Xnmos_5p04310591302098_3v512x8m81_0 pmos_5p04310591302095_3v512x8m81_0/D ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D
+ ypass_gate_3v512x8m81_0_0/pmos_5p0431059130201_3v512x8m81_0/D ypass_gate_3v512x8m81_0_0/vss
+ ypass_gate_3v512x8m81_0_0/vss nmos_5p04310591302098_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_15 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_15/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_26 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_26/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_37 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_37/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_37/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_48 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_48/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_48/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_59 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_59/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_59/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_R_3v512x8m81_19 a_n547_48# ypass_gate_3v512x8m81_0_0/vss a_16524_2#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# ypass_gate_3v512x8m81_0_0/bb ypass_gate_3v512x8m81_0_0/b
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_16 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_16/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_27 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_27/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_38 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_38/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_38/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_49 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_49/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_49/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_17 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_17/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_28 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_28/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_39 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ 018SRAM_cell1_3v512x8m81_1/w_30_512# a_16524_38786# 018SRAM_cell1_dummy_3v512x8m81_39/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_39/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_18 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_18/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_29 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_29/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_19 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_19/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_0 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_0/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_3v512x8m81_0 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ a_n547_48# 018SRAM_cell1_3v512x8m81_0/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_3v512x8m81_1/a_110_96# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_1 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_1/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_3v512x8m81_1 a_16524_38786# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_1/w_30_512#
+ a_n547_1214# 018SRAM_cell1_3v512x8m81_1/w_30_512# 018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_3v512x8m81_1/a_110_96# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_3v512x8m81
Xpmos_5p04310591302097_3v512x8m81_0 pmos_5p04310591302097_3v512x8m81_0/D pmos_5p04310591302095_3v512x8m81_0/D
+ pmos_5p04310591302095_3v512x8m81_0/D w_15880_n13729# pmos_5p04310591302097_3v512x8m81_0/S
+ pmos_5p04310591302097_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_2 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_2/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_3 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_3/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_4 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_4/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
X018SRAM_cell1_dummy_3v512x8m81_5 a_n547_48# ypass_gate_3v512x8m81_0_0/vss 018SRAM_cell1_3v512x8m81_0/w_30_512#
+ 018SRAM_cell1_3v512x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v512x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v512x8m81_5/m2_134_89# ypass_gate_3v512x8m81_0_0/vss x018SRAM_cell1_dummy_3v512x8m81
.ends

.subckt rarray4_512_3v512x8m81 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_20401#
+ m3_n1397_33733# 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96# m3_n1397_19189#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96# m3_n1397_18475#
+ m3_n1397_9493# 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_15553# 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_11917# m3_n1397_34945# 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_5143# 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_26959# 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_22111# 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_4645# m3_n1397_3931# 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_38581#
+ m3_n1397_34231# 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_16765# 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_3433# 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96# m3_n1397_19687#
+ m3_n1397_30097# 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_27673#
+ m3_n1397_36655# m3_n1397_33019# m3_n1397_7069# m3_n1397_25747# 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_247# m3_n1397_12415# 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_24037# 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_2221# 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_31309# m3_n1397_23323# m3_n1397_28171# m3_n1397_14839# 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_31807# 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_2719# m3_n1397_5857# 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_21613#
+ m3_n1397_22825# 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_1009# 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_13129# m3_n1397_17977# 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_8281# m3_n1397_1507# 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_29383# m3_n1397_8779# m3_n1397_37369# 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_37867# m3_n1397_35443# m3_n1397_9991# 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_26461# 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_28885# 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_11203#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# m3_n1397_6355#
+ m3_n1397_7567# m3_n1397_17263# m3_n1397_14341# m3_n1397_32521# 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ m3_n1397_16051# m3_n1397_25249# m3_n1397_36157# 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# m3_n1397_24535# m3_n1397_20899#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96# 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96#
+ m3_n1397_30595# VSUBS
X018SRAM_cell1_2x_3v512x8m81_608 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_619 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_427 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_405 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_438 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_449 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_416 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_983 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_961 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_950 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_972 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_994 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_235 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_202 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_213 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_224 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_268 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_246 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_279 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_257 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_780 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_791 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_609 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_90 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_428 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_406 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_417 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_439 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_940 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_984 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_962 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_951 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_973 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_995 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_203 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_236 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_225 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_214 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_247 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_269 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_258 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_770 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_792 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_781 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_91 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_80 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_407 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_429 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_418 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_941 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_985 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_930 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_963 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_952 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_974 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_996 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_204 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_226 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_237 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_215 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_248 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_259 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_760 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_782 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_771 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_793 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_590 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_92 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_81 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_70 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_408 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_419 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_920 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_942 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_986 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_931 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_953 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_975 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_997 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_964 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_216 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_205 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_227 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_238 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_249 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_761 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_750 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_783 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_772 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_794 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_580 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_591 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_93 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_71 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_82 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_60 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_409 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_921 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_910 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_943 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_987 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_954 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_932 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_976 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_998 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_965 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_217 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_206 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_239 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_228 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_762 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_751 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_740 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_784 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_795 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_773 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_581 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_592 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_570 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_50 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_94 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_83 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_72 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_61 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_900 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_922 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_944 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_988 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_911 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_955 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_933 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_977 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_999 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_966 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_207 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_229 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_218 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_763 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_752 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_730 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_741 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_785 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_796 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_774 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_560 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_582 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_593 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_571 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_390 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_40 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_51 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_95 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_84 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_73 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_62 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_901 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_934 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_923 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_945 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_989 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_912 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_956 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_978 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_967 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_208 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_764 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_753 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_731 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_742 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_720 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_219 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_786 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_797 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_775 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_561 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_583 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_550 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_572 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_594 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_391 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_380 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_41 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_52 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_30 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_96 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_85 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_74 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_63 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_902 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_935 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_924 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_946 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_913 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_957 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_979 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_968 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_209 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_765 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_743 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_721 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_754 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_732 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_798 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_787 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_776 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_710 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_562 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_584 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_540 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_551 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_573 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_595 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_392 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_370 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_381 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_0 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_42 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_53 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_20 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_31 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_97 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_86 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_75 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_64 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_903 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_936 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_925 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_947 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_914 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_958 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_969 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_766 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_744 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_755 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_733 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_722 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_799 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_777 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_788 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_700 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_711 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_552 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_530 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_541 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_563 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_585 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_574 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_596 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_393 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_371 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_360 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_382 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_190 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_43 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_10 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_54 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_21 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_32 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_76 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_98 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_87 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_65 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_904 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_937 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_926 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_915 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_948 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_959 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_745 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_767 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_756 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_734 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_723 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_789 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_778 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_712 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_701 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_520 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_553 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_531 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_542 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_586 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_564 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_575 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_597 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_372 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_350 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_394 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_361 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_383 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_2 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_191 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_180 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_44 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_11 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_55 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_22 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_33 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_77 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_66 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_88 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_99 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_927 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_905 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_916 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_949 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_938 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_746 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_724 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_757 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_735 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_768 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_779 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_702 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_713 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_510 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_532 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_543 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_587 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_565 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_576 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_598 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_554 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_521 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1020 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_351 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_395 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_362 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_340 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_384 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_373 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_3 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_192 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_181 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_170 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_45 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_12 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_34 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_23 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_56 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_89 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_78 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_67 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_906 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_917 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_928 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_939 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_725 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_758 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_736 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_747 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_769 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_703 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_714 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_522 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_511 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_599 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_555 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_533 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_544 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_588 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_566 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_577 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_500 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1010 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1021 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_374 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_352 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_396 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_341 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_330 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_363 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_385 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_4 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_160 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_171 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_193 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_182 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_46 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_13 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_35 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_24 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_79 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_68 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_57 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_907 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_918 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_929 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_737 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_759 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_748 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_726 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_704 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_715 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_501 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_523 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_512 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_556 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_534 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_578 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_589 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_545 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_567 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1011 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1000 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1022 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_375 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_320 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_353 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_397 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_386 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_364 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_342 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_331 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_5 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_194 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_183 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_161 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_172 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_150 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_14 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_47 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_36 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_25 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_69 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_58 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_919 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_908 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_727 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_749 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_738 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_705 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_716 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_502 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_513 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_535 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_524 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_557 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_546 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_579 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_568 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1012 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1023 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_376 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_310 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_354 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_398 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_387 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_365 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1001 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_343 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_321 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_332 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_6 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_184 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_195 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_162 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_173 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_140 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_151 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_15 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_48 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_37 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_26 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_59 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_909 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_728 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_739 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_706 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_717 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_503 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_514 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_558 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_536 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_547 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_569 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_525 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1013 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_377 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_311 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_344 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_399 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_300 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_333 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_388 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_366 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1002 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_322 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_355 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_7 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_196 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_185 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_163 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_174 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_130 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_141 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_152 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_49 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_38 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_27 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_16 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_729 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_707 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_718 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_504 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_515 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_559 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_537 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_548 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_526 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1014 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_301 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1003 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_345 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_334 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_389 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_378 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_367 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_323 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_312 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_356 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_8 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_890 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_197 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_186 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_164 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_175 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_131 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_142 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_153 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_120 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_39 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_17 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_28 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_708 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_719 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_505 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_516 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_538 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_549 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_527 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1015 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1004 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_346 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_379 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_302 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_335 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_368 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_324 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_313 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_357 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_891 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_880 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_9 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_165 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_176 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_132 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_154 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_110 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_121 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_143 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_198 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_187 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_18 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_29 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_709 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_506 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_517 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_539 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_528 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1016 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1005 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_347 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_303 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_336 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_369 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_325 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_314 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_358 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_892 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_881 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_870 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_188 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_199 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_166 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_177 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_155 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_122 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_133 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_100 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_111 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_144 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_19 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_518 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_507 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_529 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1017 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_326 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1006 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_348 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_304 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_337 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_315 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_359 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_893 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_882 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_860 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_871 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_167 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_189 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_178 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_112 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_134 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_123 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_101 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_145 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_156 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_690 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_519 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_508 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1018 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1007 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_349 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_327 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_305 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_338 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_316 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_894 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_872 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_883 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_861 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_850 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_168 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_179 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_33/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_124 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_102 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_146 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_113 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_157 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_135 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_680 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_691 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_509 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1008 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1019 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_306 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_317 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_873 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_862 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_851 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_840 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_328 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_339 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_895 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_884 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_169 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_114 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_125 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_103 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_147 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_136 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_158 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_670 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_681 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_692 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_1009 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_307 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_329 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_318 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_896 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_874 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_885 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_830 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_863 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_852 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_841 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_115 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_137 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_126 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_104 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_148 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_159 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_671 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_660 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_682 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_693 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_490 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_308 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_319 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_897 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_875 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_886 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_831 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_864 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_820 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_853 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_842 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_116 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_138 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_105 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_149 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_127 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_672 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_661 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_683 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_694 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_650 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_491 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_480 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_309 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_898 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_876 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_887 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_843 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_832 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_810 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_865 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_821 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_854 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_139 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_117 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_128 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_106 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_673 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_684 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_662 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_695 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_651 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_640 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_492 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_481 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_470 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_899 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_877 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_888 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_833 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_866 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_822 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_811 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_800 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_855 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_844 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_118 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_129 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_107 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_674 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_685 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_663 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_696 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_630 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_652 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_641 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_493 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_482 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_471 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_460 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_290 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_878 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_834 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_823 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_812 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_867 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_856 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_845 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_801 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_889 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_119 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_108 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_664 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_675 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_697 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_686 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_620 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_631 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_653 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_642 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_483 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_494 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_472 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_461 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_450 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_280 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_291 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_879 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_835 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_96/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_824 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_857 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_868 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_846 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_813 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_802 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_109 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_665 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_676 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_698 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_632 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_687 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_643 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_621 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_610 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_654 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_473 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_462 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_484 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_440 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_495 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_451 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_270 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_281 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_292 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_825 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_869 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_858 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_847 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_836 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_814 m3_n1397_26959# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26959# m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_27673# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_803 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_633 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_600 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_611 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_622 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_644 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_655 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_666 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_699 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_677 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_688 m3_n1397_28171# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28171# m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_28885# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_474 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_485 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_441 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_463 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_430 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_452 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_496 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_271 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_293 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_260 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_282 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_815 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_848 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_804 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_859 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_826 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_837 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_656 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_645 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_667 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_678 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_634 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_601 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_612 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_689 m3_n1397_29383# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_29383# m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30097# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_623 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_486 m3_n1397_22111# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22111# m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_22825# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_442 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_431 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_420 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_475 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_719/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_464 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_453 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_497 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_272 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_294 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_250 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_261 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_283 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_849 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_805 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_827 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_838 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_816 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_646 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_668 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_657 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_679 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_635 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_602 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_624 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_613 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_410 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_487 m3_n1397_23323# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_23323# m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24037# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_432 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_443 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_465 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_476 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_454 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_421 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_498 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_273 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_240 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_295 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_251 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_262 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_284 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_806 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_828 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_839 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_817 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_647 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_669 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_658 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_636 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_625 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_603 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_614 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_488 m3_n1397_24535# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_24535# m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25249# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_400 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_444 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_433 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_466 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_477 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_715/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_455 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_422 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_499 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_411 m3_n1397_11203# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11203# m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_230 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_274 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_241 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_252 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_296 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_263 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_285 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_807 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_81/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_829 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_818 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_82/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_637 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_659 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_626 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_604 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_615 m3_n1397_33019# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33019# m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_33733# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_648 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_489 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_401 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_478 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_445 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_434 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_456 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_467 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_423 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_412 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_990 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_220 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_231 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_264 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_242 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_275 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_253 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_297 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_286 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_819 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_89/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_808 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_99/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_605 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_627 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_616 m3_n1397_34231# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34231# m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_34945# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_649 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_638 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_402 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_479 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_446 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_435 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_468 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_457 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_424 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_413 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_980 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_991 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_221 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_210 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_232 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_265 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_243 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_276 m3_n1397_247# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_247# m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# VSUBS
+ m3_n1397_1009# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_254 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_298 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_287 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_809 m3_n1397_20899# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20899# m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_21613# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_606 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_628 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_713/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_617 m3_n1397_35443# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_35443# m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36157# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_639 m3_n1397_31807# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31807# m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_32521# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_403 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_436 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_458 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_447 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_469 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_425 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_414 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_981 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_8/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_970 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_992 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_200 m3_n1397_13627# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13627# m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_222 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_211 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_9/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_233 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_65/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_266 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_244 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_277 m3_n1397_2719# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2719# m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_973/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_255 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_299 m3_n1397_3931# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_3931# m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_288 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_607 m3_n1397_37867# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37867# m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_38581# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_717/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_629 m3_n1397_30595# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_30595# m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_31309# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_997/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_618 m3_n1397_36655# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_36655# m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_37369# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_999/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_404 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_979/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_426 m3_n1397_17263# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17263# m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_967/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_415 m3_n1397_16051# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16051# m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_965/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_982 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_46/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_960 m3_n1397_18475# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_18475# m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_6/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_971 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_459 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_437 m3_n1397_12415# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_12415# m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_448 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_995/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_993 m3_n1397_19687# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_19687# m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_20401# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_993/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_201 m3_n1397_14839# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_14839# m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_55/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_234 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_49/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_223 m3_n1397_9991# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9991# m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_23/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_212 m3_n1397_8779# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8779# m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_98/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_267 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_977/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_245 m3_n1397_6355# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_6355# m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_969/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_289 m3_n1397_5143# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5143# m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_278 m3_n1397_1507# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_1507# m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_971/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_256 m3_n1397_7567# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_7567# m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_975/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
X018SRAM_cell1_2x_3v512x8m81_790 m3_n1397_25747# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_25747# m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ VSUBS m3_n1397_26461# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512# 018SRAM_strap1_bndry_3v512x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_430_96# VSUBS 018SRAM_cell1_2x_3v512x8m81_62/018SRAM_cell1_3v512x8m81_1/a_110_96#
+ x018SRAM_cell1_2x_3v512x8m81
.ends

.subckt rcol4_512_3v512x8m81 WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[42] WL[48]
+ WL[50] WL[52] WL[54] WL[56] WL[51] WL[29] WL[20] WL[27] WL[30] WL[18] WL[41] WL[15]
+ WL[38] WL[45] WL[43] WL[40] WL[39] WL[31] WL[14] WL[16] WL[26] WL[19] WL[58] WL[60]
+ WL[62] WL[28] WL[49] WL[53] WL[55] WL[12] WL[7] WL[8] WL[5] WL[10] WL[13] WL[6]
+ tblhl GWE WL[11] din[7] q[5] q[6] q[7] din[5] din[6] q[4] pcb[7] pcb[4] WEN[4] WEN[7]
+ pcb[5] WEN[5] WEN[6] saout_R_m2_3v512x8m81_1/datain saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ rarray4_512_3v512x8m81_0/m3_n1397_13129# rarray4_512_3v512x8m81_0/m3_n1397_9493#
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass saout_m2_3v512x8m81_3/din_3v512x8m81_0/men
+ rarray4_512_3v512x8m81_0/m3_n1397_11917# rarray4_512_3v512x8m81_0/m3_n1397_5143#
+ WL[57] rdummy_3v512x4_3v512x8m81_0/a_16524_2# rdummy_3v512x4_3v512x8m81_0/ypass_gate_3v512x8m81_0_0/pcb
+ rarray4_512_3v512x8m81_0/m3_n1397_35443# saout_m2_3v512x8m81_2/q rarray4_512_3v512x8m81_0/m3_n1397_3931#
+ rarray4_512_3v512x8m81_0/m3_n1397_26461# saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ WL[1] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass rarray4_512_3v512x8m81_0/m3_n1397_22111#
+ WL[21] rarray4_512_3v512x8m81_0/m3_n1397_6355# WL[59] WL[44] rarray4_512_3v512x8m81_0/m3_n1397_19687#
+ rarray4_512_3v512x8m81_0/m3_n1397_36655# WL[9] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ rarray4_512_3v512x8m81_0/m3_n1397_27673# WL[2] rarray4_512_3v512x8m81_0/m3_n1397_24037#
+ rarray4_512_3v512x8m81_0/m3_n1397_23323# WL[0] WL[23] WL[22] rdummy_3v512x4_3v512x8m81_0/a_16524_38786#
+ rarray4_512_3v512x8m81_0/m3_n1397_7567# saout_R_m2_3v512x8m81_3/datain saout_m2_3v512x8m81_3/GWEN
+ saout_R_m2_3v512x8m81_1/sa_3v512x8m81_0/pcb WL[46] rarray4_512_3v512x8m81_0/m3_n1397_37867#
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass rarray4_512_3v512x8m81_0/m3_n1397_28885#
+ WL[4] WL[25] rarray4_512_3v512x8m81_0/m3_n1397_25249# saout_R_m2_3v512x8m81_1/q
+ saout_m2_3v512x8m81_3/q WL[3] rarray4_512_3v512x8m81_0/m3_n1397_24535# WL[24] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ saout_R_m2_3v512x8m81_3/q rarray4_512_3v512x8m81_0/m3_n1397_8779# saout_m2_3v512x8m81_3/ypass[7]
+ WL[47] rarray4_512_3v512x8m81_0/m3_n1397_8281# WL[17] rarray4_512_3v512x8m81_0/m3_n1397_20899#
+ WL[61] rarray4_512_3v512x8m81_0/m3_n1397_10705# VSS pcb[6]
Xdcap_103_novia_3v512x8m81_0[0] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[1] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[2] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[3] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[4] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[5] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[6] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[7] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[8] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[9] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[10] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[11] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[12] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[13] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[14] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[15] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[16] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[17] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[18] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[19] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[20] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[21] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[22] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[23] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[24] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[25] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[26] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[27] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[28] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[29] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[30] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[31] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[32] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[33] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[34] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xdcap_103_novia_3v512x8m81_0[35] pcb[6] VSS pcb[6] dcap_103_novia_3v512x8m81
Xsaout_m2_3v512x8m81_2 saout_m2_3v512x8m81_2/ypass[2] saout_m2_3v512x8m81_2/ypass[3]
+ saout_m2_3v512x8m81_2/ypass[4] saout_m2_3v512x8m81_2/ypass[5] saout_m2_3v512x8m81_2/ypass[6]
+ saout_m2_3v512x8m81_3/GWEN GWE saout_m2_3v512x8m81_2/bb[1] saout_m2_3v512x8m81_2/bb[3]
+ saout_m2_3v512x8m81_2/bb[4] saout_m2_3v512x8m81_2/bb[5] saout_m2_3v512x8m81_2/bb[7]
+ saout_m2_3v512x8m81_2/bb[6] saout_m2_3v512x8m81_2/b[5] saout_m2_3v512x8m81_2/b[6]
+ saout_m2_3v512x8m81_2/b[7] saout_m2_3v512x8m81_2/b[2] saout_m2_3v512x8m81_2/q saout_m2_3v512x8m81_2/pcb
+ saout_m2_3v512x8m81_2/b[1] saout_m2_3v512x8m81_2/b[3] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN[5] saout_m2_3v512x8m81_3/din_3v512x8m81_0/men saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b saout_m2_3v512x8m81_2/bb[2]
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ GWE saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass saout_m2_3v512x8m81_3/ypass[7]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ saout_m2_3v512x8m81_2/b[4] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb VSS
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass saout_m2_3v512x8m81
Xrdummy_3v512x4_3v512x8m81_0 saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_R_m2_3v512x8m81_3/bb[4] pcb[6] saout_R_m2_3v512x8m81_1/bb[5] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ rarray4_512_3v512x8m81_0/m3_n1397_36655# pcb[6] VSS WL[55] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ VSS tblhl saout_m2_3v512x8m81_3/bb[5] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass
+ pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_9493# pcb[6] VSS WL[4] WL[5] VSS pcb[6]
+ pcb[6] VSS saout_m2_3v512x8m81_2/b[3] pcb[6] saout_m2_3v512x8m81_3/b[1] rarray4_512_3v512x8m81_0/m3_n1397_13129#
+ pcb[6] saout_m2_3v512x8m81_2/bb[3] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ VSS rarray4_512_3v512x8m81_0/m3_n1397_27673# rarray4_512_3v512x8m81_0/m3_n1397_22111#
+ VSS VSS pcb[6] pcb[6] WL[3] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ VSS saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[22] pcb[6] WL[22] pcb[6] pcb[6] VSS pcb[6] VSS pcb[6] pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb pcb[6] pcb[6]
+ saout_R_m2_3v512x8m81_1/b[6] rarray4_512_3v512x8m81_0/m3_n1397_37867# VSS saout_R_m2_3v512x8m81_3/bb[5]
+ WL[54] VSS pcb[6] pcb[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ pcb[6] saout_m2_3v512x8m81_3/b[4] WL[57] rarray4_512_3v512x8m81_0/m3_n1397_36655#
+ pcb[6] WL[3] pcb[6] rdummy_3v512x4_3v512x8m81_0/ypass_gate_3v512x8m81_0_0/pcb VSS
+ VSS WL[2] VSS pcb[6] VSS pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_3/bb[2] pcb[6] saout_m2_3v512x8m81_2/bb[5] rarray4_512_3v512x8m81_0/m3_n1397_7567#
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b rarray4_512_3v512x8m81_0/m3_n1397_20899#
+ WL[51] VSS VSS VSS rarray4_512_3v512x8m81_0/m3_n1397_20899# VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_2/bb[5] pcb[6] pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_8779#
+ pcb[6] tblhl pcb[6] WL[26] VSS VSS pcb[6] WL[29] VSS saout_R_m2_3v512x8m81_3/b[3]
+ WL[61] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb VSS
+ WL[50] VSS pcb[6] pcb[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ rdummy_3v512x4_3v512x8m81_0/ypass_gate_3v512x8m81_0_0/b saout_m2_3v512x8m81_3/b[6]
+ rarray4_512_3v512x8m81_0/m3_n1397_26461# WL[59] pcb[6] WL[9] VSS VSS rarray4_512_3v512x8m81_0/m3_n1397_6355#
+ VSS pcb[6] VSS pcb[6] pcb[6] pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b pcb[6]
+ saout_m2_3v512x8m81_2/b[4] rarray4_512_3v512x8m81_0/m3_n1397_8281# saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[40] WL[23] VSS VSS VSS WL[34] pcb[6] VSS saout_m2_3v512x8m81_2/b[1] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ pcb[6] WL[30] pcb[6] pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_9493# VSS VSS pcb[6]
+ WL[30] VSS saout_R_m2_3v512x8m81_1/b[3] pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ pcb[6] WL[44] VSS pcb[6] WL[52] VSS WL[49] rarray4_512_3v512x8m81_0/m3_n1397_8281#
+ pcb[6] VSS WL[17] VSS VSS pcb[6] pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[50] pcb[6] VSS saout_m2_3v512x8m81_2/b[6] rarray4_512_3v512x8m81_0/m3_n1397_11917#
+ WL[19] VSS VSS rarray4_512_3v512x8m81_0/m3_n1397_24535# pcb[6] WL[34] VSS VSS pcb[6]
+ pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_6355# saout_R_m2_3v512x8m81_1/bb[4] VSS
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ WL[25] WL[42] VSS VSS WL[53] saout_R_m2_3v512x8m81_3/bb[2] VSS rarray4_512_3v512x8m81_0/m3_n1397_19687#
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b VSS WL[59]
+ rarray4_512_3v512x8m81_0/m3_n1397_10705# WL[15] VSS VSS VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b WL[51] pcb[6]
+ VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[21] VSS pcb[6] WL[17] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ VSS saout_R_m2_3v512x8m81_3/bb[7] rarray4_512_3v512x8m81_0/m3_n1397_25249# pcb[6]
+ VSS WL[36] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ VSS pcb[6] WL[11] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b pcb[6] VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_R_m2_3v512x8m81_1/bb[5] WL[26] rarray4_512_3v512x8m81_0/m3_n1397_37867# pcb[6]
+ VSS VSS pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ WL[32] pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ VSS WL[48] WL[1] WL[53] VSS VSS rarray4_512_3v512x8m81_0/m3_n1397_8779# VSS saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ VSS pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ pcb[6] saout_R_m2_3v512x8m81_3/bb[7] saout_R_m2_3v512x8m81_1/bb[7] pcb[6] pcb[6]
+ WL[29] VSS WL[46] VSS rarray4_512_3v512x8m81_0/m3_n1397_11917# saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ VSS rdummy_3v512x4_3v512x8m81_0/a_16524_38786# pcb[6] pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ rarray4_512_3v512x8m81_0/m3_n1397_13129# VSS rarray4_512_3v512x8m81_0/m3_n1397_22111#
+ VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb saout_R_m2_3v512x8m81_1/b[3]
+ saout_m2_3v512x8m81_2/b[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ rarray4_512_3v512x8m81_0/m3_n1397_35443# VSS WL[15] pcb[6] VSS VSS pcb[6] saout_R_m2_3v512x8m81_1/bb[4]
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb WL[23] pcb[6]
+ VSS VSS saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[49] rarray4_512_3v512x8m81_0/m3_n1397_28885# VSS VSS rarray4_512_3v512x8m81_0/m3_n1397_7567#
+ VSS WL[0] pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ VSS saout_m2_3v512x8m81_3/b[3] pcb[6] saout_R_m2_3v512x8m81_1/b[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ saout_m2_3v512x8m81_3/bb[3] WL[27] WL[47] VSS pcb[6] VSS saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ pcb[6] pcb[6] saout_R_m2_3v512x8m81_3/b[6] pcb[6] WL[40] WL[24] VSS VSS WL[36] pcb[6]
+ VSS saout_R_m2_3v512x8m81_1/bb[2] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b WL[52] pcb[6]
+ VSS rarray4_512_3v512x8m81_0/m3_n1397_10705# pcb[6] pcb[6] VSS saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb rdummy_3v512x4_3v512x8m81_0/a_16524_2#
+ WL[24] VSS saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ WL[61] VSS WL[0] VSS pcb[6] pcb[6] WL[1] WL[44] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ pcb[6] VSS VSS saout_m2_3v512x8m81_3/bb[5] pcb[6] pcb[6] saout_R_m2_3v512x8m81_3/bb[4]
+ pcb[6] WL[42] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ VSS pcb[6] pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_26461# VSS pcb[6] pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b saout_m2_3v512x8m81_2/b[4]
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb rarray4_512_3v512x8m81_0/m3_n1397_23323#
+ VSS pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/b[1] rarray4_512_3v512x8m81_0/m3_n1397_5143# saout_R_m2_3v512x8m81_1/bb[7]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb VSS WL[5] pcb[6]
+ pcb[6] WL[27] VSS VSS pcb[6] pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_28885# saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb VSS saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/b[4] rarray4_512_3v512x8m81_0/m3_n1397_3931# rarray4_512_3v512x8m81_0/m3_n1397_24535#
+ VSS VSS pcb[6] rdummy_3v512x4_3v512x8m81_0/ypass_gate_3v512x8m81_0_0/b saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ rarray4_512_3v512x8m81_0/m3_n1397_27673# pcb[6] VSS saout_R_m2_3v512x8m81_3/bb[5]
+ WL[25] pcb[6] VSS pcb[6] pcb[6] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_2/b[3] VSS saout_m2_3v512x8m81_2/bb[3] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[28] rarray4_512_3v512x8m81_0/m3_n1397_24037# VSS VSS pcb[6] saout_R_m2_3v512x8m81_1/bb[2]
+ saout_m2_3v512x8m81_3/bb[2] pcb[6] WL[9] VSS saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b WL[7] WL[48]
+ pcb[6] VSS WL[28] rarray4_512_3v512x8m81_0/m3_n1397_3931# pcb[6] VSS saout_m2_3v512x8m81_3/ypass[7]
+ VSS VSS pcb[6] pcb[6] saout_m2_3v512x8m81_2/b[1] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ pcb[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb WL[7]
+ saout_m2_3v512x8m81_3/b[6] WL[47] pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_19687#
+ VSS VSS VSS pcb[6] pcb[6] saout_R_m2_3v512x8m81_3/b[3] pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ rarray4_512_3v512x8m81_0/m3_n1397_24037# pcb[6] pcb[6] VSS rarray4_512_3v512x8m81_0/m3_n1397_35443#
+ pcb[6] VSS saout_m2_3v512x8m81_2/bb[2] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ saout_R_m2_3v512x8m81_3/b[6] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_25249# VSS pcb[6] WL[54] VSS saout_m2_3v512x8m81_3/b[3]
+ saout_m2_3v512x8m81_3/bb[3] WL[46] WL[11] pcb[6] VSS rarray4_512_3v512x8m81_0/m3_n1397_5143#
+ VSS WL[4] pcb[6] VSS pcb[6] VSS saout_m2_3v512x8m81_2/bb[2] pcb[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b WL[19] pcb[6]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ VSS rarray4_512_3v512x8m81_0/m3_n1397_23323# WL[55] VSS VSS VSS pcb[6] pcb[6] WL[2]
+ saout_R_m2_3v512x8m81_3/bb[2] VSS WL[21] pcb[6] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ pcb[6] pcb[6] VSS WL[32] pcb[6] VSS WL[57] VSS pcb[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ rdummy_3v512x4_3v512x8m81
Xsaout_m2_3v512x8m81_3 saout_m2_3v512x8m81_3/ypass[2] saout_m2_3v512x8m81_3/ypass[3]
+ saout_m2_3v512x8m81_3/ypass[4] saout_m2_3v512x8m81_3/ypass[5] saout_m2_3v512x8m81_3/ypass[6]
+ saout_m2_3v512x8m81_3/GWEN GWE saout_m2_3v512x8m81_3/bb[1] saout_m2_3v512x8m81_3/bb[3]
+ saout_m2_3v512x8m81_3/bb[4] saout_m2_3v512x8m81_3/bb[5] saout_m2_3v512x8m81_3/bb[7]
+ saout_m2_3v512x8m81_3/bb[6] saout_m2_3v512x8m81_3/b[5] saout_m2_3v512x8m81_3/b[6]
+ saout_m2_3v512x8m81_3/b[7] saout_m2_3v512x8m81_3/b[2] saout_m2_3v512x8m81_3/q saout_m2_3v512x8m81_3/pcb
+ saout_m2_3v512x8m81_3/b[1] saout_m2_3v512x8m81_3/b[3] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN[7] saout_m2_3v512x8m81_3/din_3v512x8m81_0/men saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b saout_m2_3v512x8m81_3/bb[2]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ GWE saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass saout_m2_3v512x8m81_3/ypass[7]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass
+ saout_m2_3v512x8m81_3/b[4] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass
+ pcb[6] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb VSS
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass saout_m2_3v512x8m81
Xrarray4_512_3v512x8m81_0 saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ saout_R_m2_3v512x8m81_3/bb[7] saout_R_m2_3v512x8m81_1/bb[2] saout_m2_3v512x8m81_3/bb[5]
+ saout_R_m2_3v512x8m81_1/bb[4] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b saout_m2_3v512x8m81_3/b[6]
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb WL[32] WL[53]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[30] saout_R_m2_3v512x8m81_3/b[6] WL[29] rarray4_512_3v512x8m81_0/m3_n1397_9493#
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b WL[24] saout_m2_3v512x8m81_2/bb[5]
+ saout_R_m2_3v512x8m81_3/bb[4] saout_R_m2_3v512x8m81_1/b[6] rarray4_512_3v512x8m81_0/m3_n1397_11917#
+ WL[55] saout_m2_3v512x8m81_3/b[4] rarray4_512_3v512x8m81_0/m3_n1397_5143# saout_m2_3v512x8m81_3/bb[2]
+ WL[42] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b rarray4_512_3v512x8m81_0/m3_n1397_22111#
+ saout_m2_3v512x8m81_3/bb[3] WL[7] rarray4_512_3v512x8m81_0/m3_n1397_3931# saout_m2_3v512x8m81_2/b[1]
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb saout_R_m2_3v512x8m81_1/bb[7]
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b WL[61] WL[54]
+ saout_R_m2_3v512x8m81_3/b[3] WL[26] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ WL[5] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b
+ rarray4_512_3v512x8m81_0/m3_n1397_19687# WL[47] saout_m2_3v512x8m81_3/b[1] saout_m2_3v512x8m81_2/bb[3]
+ rarray4_512_3v512x8m81_0/m3_n1397_27673# rarray4_512_3v512x8m81_0/m3_n1397_36655#
+ WL[52] WL[11] WL[40] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/bb
+ WL[0] WL[19] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ rarray4_512_3v512x8m81_0/m3_n1397_24037# saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b
+ WL[3] saout_R_m2_3v512x8m81_1/b[3] WL[49] rarray4_512_3v512x8m81_0/m3_n1397_23323#
+ WL[44] WL[23] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ WL[50] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb WL[4]
+ WL[9] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_2/b[4] WL[34] WL[36] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_m2_3v512x8m81_3/b[3] saout_R_m2_3v512x8m81_3/bb[2] WL[1] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ rarray4_512_3v512x8m81_0/m3_n1397_13129# WL[28] saout_m2_3v512x8m81_2/bb[2] rarray4_512_3v512x8m81_0/m3_n1397_8281#
+ WL[2] saout_R_m2_3v512x8m81_1/bb[5] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb WL[46] rarray4_512_3v512x8m81_0/m3_n1397_8779#
+ WL[59] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb rarray4_512_3v512x8m81_0/m3_n1397_37867#
+ rarray4_512_3v512x8m81_0/m3_n1397_35443# WL[15] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ rarray4_512_3v512x8m81_0/m3_n1397_26461# saout_R_m2_3v512x8m81_3/bb[5] rarray4_512_3v512x8m81_0/m3_n1397_28885#
+ saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b saout_m2_3v512x8m81_2/b[6]
+ WL[17] saout_m2_3v512x8m81_2/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb WL[21]
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ rarray4_512_3v512x8m81_0/m3_n1397_6355# rarray4_512_3v512x8m81_0/m3_n1397_7567#
+ WL[27] WL[22] WL[51] saout_m2_3v512x8m81_2/b[3] WL[25] rarray4_512_3v512x8m81_0/m3_n1397_25249#
+ WL[57] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb rarray4_512_3v512x8m81_0/m3_n1397_10705#
+ pcb[6] rarray4_512_3v512x8m81_0/m3_n1397_24535# rarray4_512_3v512x8m81_0/m3_n1397_20899#
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ WL[48] VSS rarray4_512_3v512x8m81
Xsaout_R_m2_3v512x8m81_1 saout_R_m2_3v512x8m81_1/ypass[2] saout_R_m2_3v512x8m81_1/ypass[3]
+ saout_R_m2_3v512x8m81_1/ypass[4] saout_R_m2_3v512x8m81_1/ypass[5] saout_R_m2_3v512x8m81_1/ypass[6]
+ GWE saout_m2_3v512x8m81_3/GWEN saout_R_m2_3v512x8m81_1/datain saout_R_m2_3v512x8m81_1/b[6]
+ saout_R_m2_3v512x8m81_1/b[5] saout_R_m2_3v512x8m81_1/b[4] saout_R_m2_3v512x8m81_1/b[2]
+ saout_R_m2_3v512x8m81_1/b[1] saout_R_m2_3v512x8m81_1/b[0] saout_R_m2_3v512x8m81_1/bb[6]
+ saout_R_m2_3v512x8m81_1/bb[7] saout_R_m2_3v512x8m81_1/q saout_R_m2_3v512x8m81_1/bb[4]
+ saout_R_m2_3v512x8m81_1/bb[3] saout_R_m2_3v512x8m81_1/bb[0] saout_R_m2_3v512x8m81_1/bb[1]
+ saout_R_m2_3v512x8m81_1/pcb saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b saout_R_m2_3v512x8m81_1/bb[2]
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN[4] saout_R_m2_3v512x8m81_1/sa_3v512x8m81_0/pcb saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ saout_m2_3v512x8m81_3/din_3v512x8m81_0/men saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_1/bb[5] saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ saout_m2_3v512x8m81_3/ypass[7] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb VSS saout_R_m2_3v512x8m81_1/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_R_m2_3v512x8m81_1/b[3] pcb[6] VSS saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ saout_R_m2_3v512x8m81
Xsaout_R_m2_3v512x8m81_3 saout_R_m2_3v512x8m81_3/ypass[2] saout_R_m2_3v512x8m81_3/ypass[3]
+ saout_R_m2_3v512x8m81_3/ypass[4] saout_R_m2_3v512x8m81_3/ypass[5] saout_R_m2_3v512x8m81_3/ypass[6]
+ GWE saout_m2_3v512x8m81_3/GWEN saout_R_m2_3v512x8m81_3/datain saout_R_m2_3v512x8m81_3/b[6]
+ saout_R_m2_3v512x8m81_3/b[5] saout_R_m2_3v512x8m81_3/b[4] saout_R_m2_3v512x8m81_3/b[2]
+ saout_R_m2_3v512x8m81_3/b[1] saout_R_m2_3v512x8m81_3/b[0] saout_R_m2_3v512x8m81_3/bb[6]
+ saout_R_m2_3v512x8m81_3/bb[7] saout_R_m2_3v512x8m81_3/q saout_R_m2_3v512x8m81_3/bb[4]
+ saout_R_m2_3v512x8m81_3/bb[3] saout_R_m2_3v512x8m81_3/bb[0] saout_R_m2_3v512x8m81_3/bb[1]
+ saout_R_m2_3v512x8m81_3/pcb saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/b
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/b saout_R_m2_3v512x8m81_3/bb[2]
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/b saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/b
+ WEN[6] saout_R_m2_3v512x8m81_3/sa_3v512x8m81_0/pcb saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/bb
+ saout_m2_3v512x8m81_3/din_3v512x8m81_0/men saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/ypass
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/ypass saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/pmos_5p0431059130201_3v512x8m81_0/D
+ saout_R_m2_3v512x8m81_3/bb[5] saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_7/bb
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/ypass saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_3/b
+ saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_1/ypass saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_a_3v512x8m81_0/ypass
+ saout_m2_3v512x8m81_3/ypass[7] saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_4/ypass
+ saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_6/bb VSS saout_R_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_5/bb
+ saout_R_m2_3v512x8m81_3/b[3] pcb[6] VSS saout_m2_3v512x8m81_3/mux821_3v512x8m81_0/ypass_gate_3v512x8m81_2/ypass
+ saout_R_m2_3v512x8m81
.ends

.subckt pmoscap_R270_3v512x8m81 m3_770_16# a_n126_928# a_n140_236# m3_152_0# w_n226_n219#
X0 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=1.20555p pd=6.07u as=0 ps=0 w=2.565u l=2.505u
X1 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=0.6733p pd=3.09u as=0 ps=0 w=2.565u l=2.505u
.ends

.subckt nmos_5p04310591302099_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.0746p pd=10.31u as=2.0746p ps=10.31u w=4.715u l=0.28u
.ends

.subckt nmos_1p2_02_R90_3v512x8m81 nmos_5p04310591302099_3v512x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v512x8m81_0/S VSUBS
Xnmos_5p04310591302099_3v512x8m81_0 nmos_5p04310591302099_3v512x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v512x8m81_0/S VSUBS nmos_5p04310591302099_3v512x8m81
.ends

.subckt pmoscap_L1_W2_R270_3v512x8m81 m3_307_0# m3_600_0# a_597_236# a_8_928# w_n88_n38#
+ a_8_236#
X0 a_597_236# a_8_928# a_8_236# w_n88_n38# pfet_03v3 ad=1.1286p pd=6.01u as=1.1286p ps=6.01u w=2.565u l=2.505u
.ends

.subckt nmos_5p043105913020102_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_1p2_01_R270_3v512x8m81 nmos_5p043105913020102_3v512x8m81_0/S a_n14_n33#
+ nmos_5p043105913020102_3v512x8m81_0/D VSUBS
Xnmos_5p043105913020102_3v512x8m81_0 nmos_5p043105913020102_3v512x8m81_0/D a_n14_n33#
+ nmos_5p043105913020102_3v512x8m81_0/S VSUBS nmos_5p043105913020102_3v512x8m81
.ends

.subckt pmos_5p043105913020101_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt pmos_1p2_01_R90_3v512x8m81 w_n137_n63# pmos_5p043105913020101_3v512x8m81_0/S
+ a_n14_n33# pmos_5p043105913020101_3v512x8m81_0/D
Xpmos_5p043105913020101_3v512x8m81_0 pmos_5p043105913020101_3v512x8m81_0/D a_n14_n33#
+ w_n137_n63# pmos_5p043105913020101_3v512x8m81_0/S pmos_5p043105913020101_3v512x8m81
.ends

.subckt pmos_5p043105913020104_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_1p2_02_R270_3v512x8m81 a_118_n33# a_n41_n33# pmos_5p043105913020104_3v512x8m81_0/D
+ w_n138_n63# pmos_5p043105913020104_3v512x8m81_0/S
Xpmos_5p043105913020104_3v512x8m81_0 pmos_5p043105913020104_3v512x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020104_3v512x8m81_0/S pmos_5p043105913020104_3v512x8m81
.ends

.subckt nmos_5p043105913020106_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1601p pd=1.64u as=0.1601p ps=1.64u w=0.305u l=0.28u
.ends

.subckt pmos_5p043105913020105_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.28u
.ends

.subckt nmos_5p043105913020107_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.6058p pd=2.85u as=1.0252p ps=5.54u w=2.33u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=1.0252p pd=5.54u as=0.6058p ps=2.85u w=2.33u l=0.28u
.ends

.subckt pmos_5p043105913020103_3v512x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=2.0526p pd=10.21u as=1.22455p ps=5.19u w=4.665u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=1.2129p pd=5.185u as=2.0526p ps=10.21u w=4.665u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=1.22455p pd=5.19u as=1.2129p ps=5.185u w=4.665u l=0.28u
.ends

.subckt pmos_1p2_03_R270_3v512x8m81 pmos_5p043105913020103_3v512x8m81_0/D a_n69_n138#
+ w_n138_n63# a_90_n138# pmos_5p043105913020103_3v512x8m81_0/S a_251_n138#
Xpmos_5p043105913020103_3v512x8m81_0 pmos_5p043105913020103_3v512x8m81_0/D a_251_n138#
+ pmos_5p043105913020103_3v512x8m81_0/S a_n69_n138# a_90_n138# w_n138_n63# pmos_5p043105913020103_3v512x8m81
.ends

.subckt pmos_5p043105913020108_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6669p pd=3.085u as=1.1286p ps=6.01u w=2.565u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1286p pd=6.01u as=0.6669p ps=3.085u w=2.565u l=0.28u
.ends

.subckt pmos_1p2_01_R270_3v512x8m81 pmos_5p043105913020108_3v512x8m81_0/S w_n246_n93#
+ pmos_5p043105913020108_3v512x8m81_0/D a_118_n33# a_n41_n33#
Xpmos_5p043105913020108_3v512x8m81_0 pmos_5p043105913020108_3v512x8m81_0/D a_n41_n33#
+ a_118_n33# w_n246_n93# pmos_5p043105913020108_3v512x8m81_0/S pmos_5p043105913020108_3v512x8m81
.ends

.subckt nmos_1p2_02_R270_3v512x8m81 a_n14_n33# nmos_5p04310591302044_3v512x8m81_0/S
+ nmos_5p04310591302044_3v512x8m81_0/D VSUBS
Xnmos_5p04310591302044_3v512x8m81_0 nmos_5p04310591302044_3v512x8m81_0/D a_n14_n33#
+ nmos_5p04310591302044_3v512x8m81_0/S VSUBS nmos_5p04310591302044_3v512x8m81
.ends

.subckt nmos_5p043105913020109_3v512x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_5p043105913020110_3v512x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3256p pd=2.36u as=0.3256p ps=2.36u w=0.74u l=0.28u
.ends

.subckt xdec_3v512x8m81 RWL LWL men xc xb xa m2_11898_n156# m2_9070_n156# m2_7748_n156#
+ m2_8806_n156# m2_10577_n156# m2_10840_n156# m2_7219_n156# m2_7483_n156# m2_11634_n156#
+ m2_12427_n156# m2_8277_n156# m2_8541_n156# m2_11105_n156# m2_11370_n156# m2_12163_n156#
+ m2_8012_n156# vss vdd
Xpmos_1p2_02_R270_3v512x8m81_0 pmos_5p043105913020105_3v512x8m81_3/S pmos_5p043105913020105_3v512x8m81_3/S
+ men vdd nmos_5p043105913020109_3v512x8m81_0/S pmos_1p2_02_R270_3v512x8m81
Xnmos_5p043105913020106_3v512x8m81_0 vss pmos_5p043105913020105_3v512x8m81_3/S pmos_5p043105913020110_3v512x8m81_0/S
+ vss nmos_5p043105913020106_3v512x8m81
Xpmos_5p043105913020105_3v512x8m81_1 pmos_5p043105913020105_3v512x8m81_3/S xb vdd
+ vdd pmos_5p043105913020105_3v512x8m81
Xpmos_5p043105913020105_3v512x8m81_2 vdd xa vdd pmos_5p043105913020105_3v512x8m81_3/S
+ pmos_5p043105913020105_3v512x8m81
Xpmos_5p043105913020105_3v512x8m81_3 vdd xc vdd pmos_5p043105913020105_3v512x8m81_3/S
+ pmos_5p043105913020105_3v512x8m81
Xnmos_5p043105913020107_3v512x8m81_0 LWL pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D
+ pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D vss vss nmos_5p043105913020107_3v512x8m81
Xpmos_1p2_03_R270_3v512x8m81_0 vdd pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D
+ vdd pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D LWL pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D
+ pmos_1p2_03_R270_3v512x8m81
Xnmos_5p043105913020107_3v512x8m81_1 RWL pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D
+ pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D vss vss nmos_5p043105913020107_3v512x8m81
Xpmos_1p2_01_R270_3v512x8m81_0 vdd vdd pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D
+ nmos_5p043105913020109_3v512x8m81_0/S nmos_5p043105913020109_3v512x8m81_0/S pmos_1p2_01_R270_3v512x8m81
Xpmos_1p2_01_R270_3v512x8m81_1 vdd vdd pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D
+ nmos_5p043105913020109_3v512x8m81_0/S nmos_5p043105913020109_3v512x8m81_0/S pmos_1p2_01_R270_3v512x8m81
Xnmos_1p2_02_R270_3v512x8m81_0 pmos_5p043105913020105_3v512x8m81_3/S nmos_5p043105913020109_3v512x8m81_0/S
+ vss vss nmos_1p2_02_R270_3v512x8m81
Xnmos_5p043105913020109_3v512x8m81_0 men pmos_5p043105913020110_3v512x8m81_0/S pmos_5p043105913020110_3v512x8m81_0/S
+ nmos_5p043105913020109_3v512x8m81_0/S vss nmos_5p043105913020109_3v512x8m81
Xpmos_5p043105913020103_3v512x8m81_0 vdd pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D
+ RWL pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D
+ vdd pmos_5p043105913020103_3v512x8m81
Xpmos_5p043105913020110_3v512x8m81_0 vdd pmos_5p043105913020105_3v512x8m81_3/S vdd
+ pmos_5p043105913020110_3v512x8m81_0/S pmos_5p043105913020110_3v512x8m81
X0 vss xc a_9450_422# vss nfet_03v3 ad=0.88935p pd=4.15u as=0.29032p ps=1.865u w=1.47u l=0.28u
X1 vss nmos_5p043105913020109_3v512x8m81_0/S pmos_1p2_01_R270_3v512x8m81_1/pmos_5p043105913020108_3v512x8m81_0/D vss nfet_03v3 ad=0.2796p pd=4.9u as=1.0252p ps=5.54u w=2.33u l=0.28u
X2 a_9450_280# xa pmos_5p043105913020105_3v512x8m81_3/S vss nfet_03v3 ad=0.31605p pd=1.9u as=0.74235p ps=3.95u w=1.47u l=0.28u
X3 a_9450_422# xb a_9450_280# vss nfet_03v3 ad=0.29032p pd=1.865u as=0.31605p ps=1.9u w=1.47u l=0.28u
X4 vss nmos_5p043105913020109_3v512x8m81_0/S pmos_1p2_01_R270_3v512x8m81_0/pmos_5p043105913020108_3v512x8m81_0/D vss nfet_03v3 ad=1.15335p pd=5.65u as=1.0718p ps=5.58u w=2.33u l=0.28u
.ends

.subckt xdec8_3v512x8m81 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] LWL[1] LWL[7] LWL[6]
+ LWL[0] LWL[3] xa[3] xa[6] xa[0] xa[5] xa[2] xdec_3v512x8m81_7/m2_10577_n156# RWL[3]
+ xdec_3v512x8m81_7/m2_11634_n156# RWL[0] xdec_3v512x8m81_7/m2_12427_n156# xc xdec_3v512x8m81_7/m2_8277_n156#
+ RWL[6] xdec_3v512x8m81_7/m2_8012_n156# xa[1] xb xa[7] xdec_3v512x8m81_7/m2_10840_n156#
+ xa[4] men xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_7483_n156# RWL[1] xdec_3v512x8m81_7/m2_9070_n156#
+ xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_11105_n156# vdd xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_11898_n156# RWL[7] vss
Xxdec_3v512x8m81_0 RWL[6] LWL[6] men xc xb xa[6] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_1 RWL[4] LWL[4] men xc xb xa[4] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_2 RWL[2] LWL[2] men xc xb xa[2] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_3 RWL[0] LWL[0] men xc xb xa[0] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_4 RWL[7] LWL[7] men xc xb xa[7] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_5 RWL[5] LWL[5] men xc xb xa[5] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_6 RWL[3] LWL[3] men xc xb xa[3] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
Xxdec_3v512x8m81_7 RWL[1] LWL[1] men xc xb xa[1] xdec_3v512x8m81_7/m2_11898_n156#
+ xdec_3v512x8m81_7/m2_9070_n156# xdec_3v512x8m81_7/m2_7748_n156# xdec_3v512x8m81_7/m2_8806_n156#
+ xdec_3v512x8m81_7/m2_10577_n156# xdec_3v512x8m81_7/m2_10840_n156# xdec_3v512x8m81_7/m2_7219_n156#
+ xdec_3v512x8m81_7/m2_7483_n156# xdec_3v512x8m81_7/m2_11634_n156# xdec_3v512x8m81_7/m2_12427_n156#
+ xdec_3v512x8m81_7/m2_8277_n156# xdec_3v512x8m81_7/m2_8541_n156# xdec_3v512x8m81_7/m2_11105_n156#
+ xdec_3v512x8m81_7/m2_11370_n156# xdec_3v512x8m81_7/m2_12163_n156# xdec_3v512x8m81_7/m2_8012_n156#
+ vss vdd xdec_3v512x8m81
.ends

.subckt xdec32_3v512x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[13] RWL[12] LWL[9]
+ LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[5] RWL[3] RWL[2]
+ LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6] LWL[28]
+ LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19] RWL[23]
+ RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xb[2] xb[0] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[20] RWL[24] RWL[21] RWL[0] RWL[25] xa[1] xa[3] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7748_n156#
+ xa[0] xa[2] RWL[28] RWL[8] RWL[1] xc men RWL[14] RWL[7] xb[1] RWL[4] RWL[16] xa[5]
+ RWL[29] RWL[9] xa[7] RWL[22] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156#
+ vss xa[4] xb[3] vdd xa[6]
Xxdec8_3v512x8m81_0 LWL[29] LWL[28] LWL[26] RWL[29] RWL[28] RWL[26] LWL[25] LWL[31]
+ LWL[30] LWL[24] LWL[27] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[27] xa[3] RWL[24]
+ xa[0] xc xb[3] RWL[30] xc xa[1] xb[3] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1]
+ xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156# RWL[25] xb[0] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7748_n156#
+ xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2] RWL[31] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_1 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] LWL[1] LWL[7] LWL[6]
+ LWL[0] LWL[3] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[3] xa[3] RWL[0] xa[0] xc xb[3]
+ RWL[6] xc xa[1] xb[0] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[1] xb[0] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7748_n156# xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156#
+ xa[2] RWL[7] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_2 LWL[13] LWL[12] LWL[10] RWL[13] RWL[12] RWL[10] LWL[9] LWL[15]
+ LWL[14] LWL[8] LWL[11] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[11] xa[3] RWL[8]
+ xa[0] xc xb[3] RWL[14] xc xa[1] xb[1] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1]
+ xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156# RWL[9] xb[0] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7748_n156#
+ xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2] RWL[15] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_3 LWL[21] LWL[20] LWL[18] RWL[21] RWL[20] RWL[18] LWL[17] LWL[23]
+ LWL[22] LWL[16] LWL[19] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[19] xa[3] RWL[16]
+ xa[0] xc xb[3] RWL[22] xc xa[1] xb[2] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1]
+ xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156# RWL[17] xb[0] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7748_n156#
+ xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2] RWL[23] vss xdec8_3v512x8m81
.ends

.subckt xdec32_468_3v512x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[13] RWL[12]
+ LWL[9] LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[5] RWL[3]
+ RWL[1] RWL[0] RWL[2] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11]
+ LWL[10] RWL[6] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20]
+ LWL[19] RWL[23] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19]
+ xa[2] xb[2] xb[1] xb[0] xc xa[1] RWL[20] RWL[24] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_8012_n156#
+ xa[7] RWL[21] xa[6] RWL[25] xa[3] xa[0] RWL[8] RWL[28] RWL[14] men RWL[7] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[16] RWL[4] xa[5] RWL[29] RWL[9] RWL[22] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156#
+ vss xa[4] xb[3] vdd
Xxdec8_3v512x8m81_0 LWL[29] LWL[28] LWL[26] RWL[29] RWL[28] RWL[26] LWL[25] LWL[31]
+ LWL[30] LWL[24] LWL[27] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[27] xa[3] RWL[24]
+ xa[0] xc xb[3] RWL[30] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_8012_n156# xa[1]
+ xb[3] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[25] xb[0] xc xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2]
+ RWL[31] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_1 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] LWL[1] LWL[7] LWL[6]
+ LWL[0] LWL[3] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[3] xa[3] RWL[0] xa[0] xc xb[3]
+ RWL[6] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_8012_n156# xa[1] xb[0] xa[7] xa[6]
+ xa[4] men xa[4] xb[2] xb[1] xa[1] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[1] xb[0] xc xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2]
+ RWL[7] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_2 LWL[13] LWL[12] LWL[10] RWL[13] RWL[12] RWL[10] LWL[9] LWL[15]
+ LWL[14] LWL[8] LWL[11] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[11] xa[3] RWL[8]
+ xa[0] xc xb[3] RWL[14] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_8012_n156# xa[1]
+ xb[1] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[9] xb[0] xc xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2]
+ RWL[15] vss xdec8_3v512x8m81
Xxdec8_3v512x8m81_3 LWL[21] LWL[20] LWL[18] RWL[21] RWL[20] RWL[18] LWL[17] LWL[23]
+ LWL[22] LWL[16] LWL[19] xa[3] xa[6] xa[0] xa[5] xa[2] xa[7] RWL[19] xa[3] RWL[16]
+ xa[0] xc xb[3] RWL[22] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_8012_n156# xa[1]
+ xb[2] xa[7] xa[6] xa[4] men xa[4] xb[2] xb[1] xa[1] xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7483_n156#
+ RWL[17] xb[0] xc xa[5] vdd xdec8_3v512x8m81_3/xdec_3v512x8m81_7/m2_7219_n156# xa[2]
+ RWL[23] vss xdec8_3v512x8m81
.ends

.subckt pmos_5p043105913020100_3v512x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.5314p pd=6.41u as=2.5916p ps=12.66u w=5.89u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=2.5916p pd=12.66u as=1.5314p ps=6.41u w=5.89u l=0.28u
.ends

.subckt pmos_1p2_02_R90_3v512x8m81 pmos_5p043105913020100_3v512x8m81_0/D a_118_n33#
+ a_n41_n33# pmos_5p043105913020100_3v512x8m81_0/S w_n138_n63#
Xpmos_5p043105913020100_3v512x8m81_0 pmos_5p043105913020100_3v512x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020100_3v512x8m81_0/S pmos_5p043105913020100_3v512x8m81
.ends

.subckt nmos_5p043105913020111_3v512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.5412p pd=3.34u as=0.5412p ps=3.34u w=1.23u l=0.28u
.ends

.subckt xdec64_3v512x8m81 DRWL RWL[34] RWL[35] RWL[36] RWL[37] RWL[38] RWL[39] RWL[40]
+ RWL[42] RWL[44] RWL[47] RWL[49] RWL[50] RWL[51] RWL[52] RWL[53] RWL[54] RWL[55]
+ RWL[56] RWL[57] RWL[58] RWL[60] RWL[62] LWL[62] LWL[61] LWL[57] LWL[55] LWL[53]
+ LWL[52] LWL[50] LWL[49] LWL[48] LWL[37] LWL[35] DLWL LWL[19] LWL[20] LWL[21] LWL[22]
+ LWL[26] LWL[10] LWL[12] LWL[14] LWL[15] LWL[17] LWL[18] LWL[5] LWL[4] LWL[3] LWL[8]
+ LWL[9] LWL[6] LWL[7] RWL[31] RWL[25] RWL[6] RWL[4] RWL[5] RWL[7] RWL[8] RWL[10]
+ RWL[12] RWL[13] RWL[14] RWL[15] xb[0] xb[1] xb[2] xb[3] xa[7] xa[6] xa[5] xa[4]
+ xa[0] men xa[3] xa[2] xa[1] xc[0] xc[1] LWL[24] RWL[59] LWL[45] LWL[29] LWL[63]
+ RWL[28] RWL[23] LWL[46] LWL[43] RWL[26] LWL[27] RWL[45] LWL[44] RWL[24] xdec32_468_3v512x8m81_0/LWL[29]
+ RWL[2] xdec32_468_3v512x8m81_0/LWL[30] LWL[42] LWL[33] RWL[3] LWL[13] RWL[22] RWL[11]
+ RWL[21] RWL[63] LWL[32] LWL[2] RWL[29] RWL[0] LWL[41] LWL[60] LWL[40] LWL[25] RWL[20]
+ LWL[1] RWL[43] LWL[0] RWL[32] RWL[30] LWL[58] LWL[38] LWL[51] RWL[48] RWL[18] vdd
+ LWL[59] LWL[30] RWL[33] RWL[1] LWL[56] LWL[11] LWL[36] RWL[19] RWL[9] RWL[61] RWL[46]
+ LWL[16] RWL[17] RWL[27] LWL[39] LWL[28] LWL[47] RWL[16] LWL[23] LWL[54] LWL[34]
+ vss LWL[31] RWL[41]
Xpmoscap_R270_3v512x8m81_5 RWL[6] vss vdd RWL[7] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_6 RWL[4] vss vdd RWL[5] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_7 RWL[2] vss vdd RWL[3] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_8 RWL[0] vss vdd RWL[1] vdd pmoscap_R270_3v512x8m81
Xnmos_1p2_02_R90_3v512x8m81_0 vss nmos_5p043105913020111_3v512x8m81_0/S DLWL vss nmos_1p2_02_R90_3v512x8m81
Xpmoscap_R270_3v512x8m81_50 RWL[56] vss vdd RWL[57] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_60 RWL[36] vss vdd RWL[37] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_61 RWL[34] vss vdd RWL[35] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_9 RWL[30] vss vdd RWL[31] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_51 RWL[54] vss vdd RWL[55] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_40 LWL[46] vss vdd LWL[47] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_62 LWL[32] vss vdd LWL[33] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_52 RWL[52] vss vdd RWL[53] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_41 LWL[44] vss vdd LWL[45] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_63 RWL[32] vss vdd RWL[33] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_30 LWL[20] vss vdd LWL[21] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_53 RWL[50] vss vdd RWL[51] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_42 LWL[42] vss vdd LWL[43] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_31 LWL[18] vss vdd LWL[19] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_20 LWL[8] vss vdd LWL[9] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_32 xdec32_468_3v512x8m81_0/LWL[30] vss vdd LWL[63] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_54 RWL[48] vss vdd RWL[49] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_43 LWL[40] vss vdd LWL[41] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_10 RWL[28] vss vdd RWL[29] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_21 LWL[6] vss vdd LWL[7] vdd pmoscap_R270_3v512x8m81
Xpmoscap_L1_W2_R270_3v512x8m81_0 DLWL vdd vdd vss vdd vdd pmoscap_L1_W2_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_33 LWL[60] vss vdd xdec32_468_3v512x8m81_0/LWL[29] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_55 RWL[46] vss vdd RWL[47] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_44 LWL[38] vss vdd LWL[39] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_11 RWL[26] vss vdd RWL[27] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_22 LWL[4] vss vdd LWL[5] vdd pmoscap_R270_3v512x8m81
Xpmoscap_L1_W2_R270_3v512x8m81_1 DRWL vdd vdd vss vdd vdd pmoscap_L1_W2_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_34 LWL[58] vss vdd LWL[59] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_56 RWL[44] vss vdd RWL[45] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_45 LWL[36] vss vdd LWL[37] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_12 RWL[24] vss vdd RWL[25] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_23 LWL[2] vss vdd LWL[3] vdd pmoscap_R270_3v512x8m81
Xnmos_1p2_01_R270_3v512x8m81_0 pmos_5p043105913020101_3v512x8m81_1/D vdd men vss nmos_1p2_01_R270_3v512x8m81
Xpmos_1p2_01_R90_3v512x8m81_0 vdd nmos_5p043105913020111_3v512x8m81_0/S pmos_5p043105913020101_3v512x8m81_1/D
+ vdd pmos_1p2_01_R90_3v512x8m81
Xpmoscap_R270_3v512x8m81_35 LWL[56] vss vdd LWL[57] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_57 RWL[42] vss vdd RWL[43] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_46 LWL[34] vss vdd LWL[35] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_13 RWL[22] vss vdd RWL[23] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_24 LWL[0] vss vdd LWL[1] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_47 RWL[62] vss vdd RWL[63] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_48 RWL[60] vss vdd RWL[61] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_36 LWL[54] vss vdd LWL[55] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_37 LWL[52] vss vdd LWL[53] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_58 RWL[40] vss vdd RWL[41] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_59 RWL[38] vss vdd RWL[39] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_26 LWL[28] vss vdd LWL[29] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_25 LWL[30] vss vdd LWL[31] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_15 RWL[18] vss vdd RWL[19] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_14 RWL[20] vss vdd RWL[21] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_49 RWL[58] vss vdd RWL[59] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_38 LWL[50] vss vdd LWL[51] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_27 LWL[26] vss vdd LWL[27] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_16 LWL[16] vss vdd LWL[17] vdd pmoscap_R270_3v512x8m81
Xpmos_5p043105913020101_3v512x8m81_0 vdd pmos_5p043105913020101_3v512x8m81_1/D vdd
+ pmos_5p043105913020101_3v512x8m81_0/S pmos_5p043105913020101_3v512x8m81
Xpmoscap_R270_3v512x8m81_39 LWL[48] vss vdd LWL[49] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_28 LWL[24] vss vdd LWL[25] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_17 LWL[14] vss vdd LWL[15] vdd pmoscap_R270_3v512x8m81
Xpmos_5p043105913020101_3v512x8m81_1 pmos_5p043105913020101_3v512x8m81_1/D vss vdd
+ men pmos_5p043105913020101_3v512x8m81
Xpmoscap_R270_3v512x8m81_29 LWL[22] vss vdd LWL[23] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_18 LWL[12] vss vdd LWL[13] vdd pmoscap_R270_3v512x8m81
Xxdec32_3v512x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[13] RWL[12] LWL[9]
+ LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[5] RWL[3] RWL[2]
+ LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6] LWL[28]
+ LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19] RWL[23]
+ RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xb[2] xb[0] vdd
+ RWL[20] RWL[24] RWL[21] RWL[0] RWL[25] xa[1] xa[3] xc[1] xa[0] xa[2] RWL[28] RWL[8]
+ RWL[1] xc[0] men RWL[14] RWL[7] xb[1] RWL[4] RWL[16] xa[5] RWL[29] RWL[9] xa[7]
+ RWL[22] vdd vss xa[4] xb[3] vdd xa[6] xdec32_3v512x8m81
Xpmoscap_R270_3v512x8m81_19 LWL[10] vss vdd LWL[11] vdd pmoscap_R270_3v512x8m81
Xxdec32_468_3v512x8m81_0 LWL[38] LWL[39] RWL[50] RWL[49] RWL[47] RWL[45] RWL[44] LWL[41]
+ LWL[40] LWL[32] LWL[33] LWL[34] LWL[35] LWL[36] LWL[37] RWL[43] RWL[42] RWL[37]
+ RWL[35] RWL[33] RWL[32] RWL[34] LWL[50] LWL[49] LWL[48] LWL[47] LWL[46] LWL[45]
+ LWL[44] LWL[43] LWL[42] RWL[38] LWL[60] LWL[59] LWL[58] LWL[57] LWL[56] LWL[55]
+ LWL[54] LWL[53] LWL[52] LWL[51] RWL[55] RWL[58] RWL[59] RWL[62] RWL[63] LWL[63]
+ xdec32_468_3v512x8m81_0/LWL[30] xdec32_468_3v512x8m81_0/LWL[29] RWL[51] xa[2] xb[2]
+ xb[1] xb[0] xc[1] xa[1] RWL[52] RWL[56] xc[0] xa[7] RWL[53] xa[6] RWL[57] xa[3]
+ xa[0] RWL[40] RWL[60] RWL[46] men RWL[39] vdd RWL[48] RWL[36] xa[5] RWL[61] RWL[41]
+ RWL[54] vdd vss xa[4] xb[3] vdd xdec32_468_3v512x8m81
Xpmos_1p2_02_R90_3v512x8m81_0 DLWL nmos_5p043105913020111_3v512x8m81_0/S nmos_5p043105913020111_3v512x8m81_0/S
+ vdd vdd pmos_1p2_02_R90_3v512x8m81
Xpmos_1p2_02_R90_3v512x8m81_1 DRWL pmos_5p043105913020101_3v512x8m81_0/S pmos_5p043105913020101_3v512x8m81_0/S
+ vdd vdd pmos_1p2_02_R90_3v512x8m81
Xnmos_5p04310591302099_3v512x8m81_0 vss pmos_5p043105913020101_3v512x8m81_0/S DRWL
+ vss nmos_5p04310591302099_3v512x8m81
Xnmos_5p043105913020111_3v512x8m81_0 vss pmos_5p043105913020101_3v512x8m81_1/D nmos_5p043105913020111_3v512x8m81_0/S
+ vss nmos_5p043105913020111_3v512x8m81
Xnmos_5p043105913020111_3v512x8m81_1 vss pmos_5p043105913020101_3v512x8m81_1/D pmos_5p043105913020101_3v512x8m81_0/S
+ vss nmos_5p043105913020111_3v512x8m81
Xpmoscap_R270_3v512x8m81_0 RWL[16] vss vdd RWL[17] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_1 RWL[14] vss vdd RWL[15] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_2 RWL[12] vss vdd RWL[13] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_3 RWL[10] vss vdd RWL[11] vdd pmoscap_R270_3v512x8m81
Xpmoscap_R270_3v512x8m81_4 RWL[8] vss vdd RWL[9] vdd pmoscap_R270_3v512x8m81
.ends

.subckt gf180mcu_ocd_ip_sram__sram512x8m8wm1 GWEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1]
+ VDD WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] A[0] D[1] A[1] A[2] D[3] A[3] A[4] D[5] A[5]
+ A[6] D[7] A[7] A[8] CEN VSS WEN[0] CLK WEN[1] WEN[2] Q[0]
Xcontrol_3v512x8_3v512x8m81_0 control_3v512x8_3v512x8m81_0/RYS[7] control_3v512x8_3v512x8m81_0/RYS[6]
+ control_3v512x8_3v512x8m81_0/RYS[5] control_3v512x8_3v512x8m81_0/RYS[4] control_3v512x8_3v512x8m81_0/RYS[3]
+ control_3v512x8_3v512x8m81_0/RYS[2] control_3v512x8_3v512x8m81_0/RYS[1] control_3v512x8_3v512x8m81_0/RYS[0]
+ VSS control_3v512x8_3v512x8m81_0/LYS[1] control_3v512x8_3v512x8m81_0/LYS[2] control_3v512x8_3v512x8m81_0/LYS[3]
+ control_3v512x8_3v512x8m81_0/LYS[6] control_3v512x8_3v512x8m81_0/LYS[5] control_3v512x8_3v512x8m81_0/LYS[4]
+ control_3v512x8_3v512x8m81_0/LYS[7] rcol4_512_3v512x8m81_0/tblhl control_3v512x8_3v512x8m81_0/IGWEN
+ xdec64_3v512x8m81_0/xb[3] xdec64_3v512x8m81_0/xb[2] xdec64_3v512x8m81_0/xb[0] xdec64_3v512x8m81_0/xa[7]
+ xdec64_3v512x8m81_0/xa[6] xdec64_3v512x8m81_0/xa[5] xdec64_3v512x8m81_0/xa[4] xdec64_3v512x8m81_0/xa[3]
+ xdec64_3v512x8m81_0/xa[2] A[0] CEN xdec64_3v512x8m81_0/xb[1] control_3v512x8_3v512x8m81_0/xc[3]
+ xdec64_3v512x8m81_0/xc[1] control_3v512x8_3v512x8m81_0/xc[2] xdec64_3v512x8m81_0/xa[1]
+ VSS A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWEN lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[1]
+ lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[2] lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[4]
+ lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[5] lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[6]
+ rcol4_512_3v512x8m81_0/GWE lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[7]
+ xdec64_3v512x8m81_0/xa[0] VDD xdec64_3v512x8m81_0/xc[0] xdec64_3v512x8m81_0/men
+ VSS VDD control_3v512x8_3v512x8m81
Xlcol4_512_3v512x8m81_0 xdec64_3v512x8m81_0/LWL[33] lcol4_512_3v512x8m81_0/WL[33]
+ xdec64_3v512x8m81_0/LWL[35] lcol4_512_3v512x8m81_0/WL[38] VSS VSS xdec64_3v512x8m81_0/LWL[37]
+ VSS xdec64_3v512x8m81_0/LWL[42] VSS xdec64_3v512x8m81_0/LWL[44] lcol4_512_3v512x8m81_0/WL[43]
+ xdec64_3v512x8m81_0/LWL[46] lcol4_512_3v512x8m81_0/WL[45] xdec64_3v512x8m81_0/LWL[48]
+ xdec64_3v512x8m81_0/LWL[49] xdec64_3v512x8m81_0/LWL[52] xdec64_3v512x8m81_0/LWL[53]
+ xdec64_3v512x8m81_0/LWL[54] xdec64_3v512x8m81_0/LWL[55] xdec64_3v512x8m81_0/LWL[56]
+ xdec64_3v512x8m81_0/LWL[57] lcol4_512_3v512x8m81_0/WL[56] lcol4_512_3v512x8m81_0/WL[58]
+ VSS xdec64_3v512x8m81_0/LWL[63] VSS VDD xdec64_3v512x8m81_0/LWL[26] xdec64_3v512x8m81_0/LWL[25]
+ xdec64_3v512x8m81_0/LWL[24] xdec64_3v512x8m81_0/LWL[23] xdec64_3v512x8m81_0/LWL[22]
+ lcol4_512_3v512x8m81_0/WL[20] lcol4_512_3v512x8m81_0/WL[18] xdec64_3v512x8m81_0/LWL[18]
+ VSS xdec64_3v512x8m81_0/LWL[16] VSS lcol4_512_3v512x8m81_0/WL[13] VSS xdec64_3v512x8m81_0/LWL[11]
+ VSS lcol4_512_3v512x8m81_0/WL[8] lcol4_512_3v512x8m81_0/WL[6] lcol4_512_3v512x8m81_0/WL[31]
+ xdec64_3v512x8m81_0/LWL[31] xdec64_3v512x8m81_0/LWL[29] xdec64_3v512x8m81_0/LWL[28]
+ xdec64_3v512x8m81_0/LWL[27] lcol4_512_3v512x8m81_0/din[1] lcol4_512_3v512x8m81_0/din[3]
+ lcol4_512_3v512x8m81_0/din[2] lcol4_512_3v512x8m81_0/q[1] lcol4_512_3v512x8m81_0/q[2]
+ lcol4_512_3v512x8m81_0/q[3] lcol4_512_3v512x8m81_0/pcb[2] lcol4_512_3v512x8m81_0/pcb[3]
+ lcol4_512_3v512x8m81_0/pcb[0] lcol4_512_3v512x8m81_0/pcb[1] WEN[0] WEN[1] WEN[2]
+ WEN[3] Q[3] xdec64_3v512x8m81_0/LWL[40] xdec64_3v512x8m81_0/LWL[41] D[3] xdec64_3v512x8m81_0/LWL[43]
+ xdec64_3v512x8m81_0/LWL[60] lcol4_512_3v512x8m81_0/WL[59] xdec64_3v512x8m81_0/LWL[45]
+ xdec64_3v512x8m81_0/xdec32_468_3v512x8m81_0/LWL[30] rcol4_512_3v512x8m81_0/GWE xdec64_3v512x8m81_0/LWL[47]
+ rcol4_512_3v512x8m81_0/GWE control_3v512x8_3v512x8m81_0/IGWEN rcol4_512_3v512x8m81_0/GWE
+ Q[2] xdec64_3v512x8m81_0/LWL[0] xdec64_3v512x8m81_0/LWL[10] xdec64_3v512x8m81_0/men
+ xdec64_3v512x8m81_0/LWL[1] xdec64_3v512x8m81_0/LWL[2] xdec64_3v512x8m81_0/LWL[12]
+ xdec64_3v512x8m81_0/LWL[3] xdec64_3v512x8m81_0/LWL[13] xdec64_3v512x8m81_0/LWL[30]
+ xdec64_3v512x8m81_0/LWL[4] xdec64_3v512x8m81_0/LWL[14] Q[1] xdec64_3v512x8m81_0/LWL[5]
+ xdec64_3v512x8m81_0/LWL[15] xdec64_3v512x8m81_0/LWL[32] xdec64_3v512x8m81_0/LWL[6]
+ xdec64_3v512x8m81_0/LWL[50] rcol4_512_3v512x8m81_0/GWE xdec64_3v512x8m81_0/LWL[7]
+ xdec64_3v512x8m81_0/LWL[17] xdec64_3v512x8m81_0/LWL[34] control_3v512x8_3v512x8m81_0/LYS[7]
+ xdec64_3v512x8m81_0/LWL[51] xdec64_3v512x8m81_0/LWL[8] lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[1]
+ xdec64_3v512x8m81_0/LWL[9] xdec64_3v512x8m81_0/LWL[19] xdec64_3v512x8m81_0/LWL[36]
+ lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[2] VDD xdec64_3v512x8m81_0/LWL[38]
+ lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[4] xdec64_3v512x8m81_0/LWL[39]
+ lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[5] lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[6]
+ Q[0] lcol4_512_3v512x8m81_0/col_512a_3v512x8m81_0/ypass[7] xdec64_3v512x8m81_0/LWL[58]
+ xdec64_3v512x8m81_0/LWL[59] rcol4_512_3v512x8m81_0/GWE D[1] xdec64_3v512x8m81_0/LWL[20]
+ VDD VSS xdec64_3v512x8m81_0/LWL[21] lcol4_512_3v512x8m81
Xrcol4_512_3v512x8m81_0 xdec64_3v512x8m81_0/RWL[33] rcol4_512_3v512x8m81_0/WL[33]
+ xdec64_3v512x8m81_0/RWL[35] rcol4_512_3v512x8m81_0/WL[35] xdec64_3v512x8m81_0/RWL[37]
+ VSS xdec64_3v512x8m81_0/RWL[44] xdec64_3v512x8m81_0/RWL[50] xdec64_3v512x8m81_0/RWL[52]
+ xdec64_3v512x8m81_0/RWL[54] xdec64_3v512x8m81_0/RWL[56] rcol4_512_3v512x8m81_0/WL[56]
+ xdec64_3v512x8m81_0/RWL[53] xdec64_3v512x8m81_0/RWL[30] rcol4_512_3v512x8m81_0/WL[20]
+ xdec64_3v512x8m81_0/RWL[28] xdec64_3v512x8m81_0/RWL[31] VSS VSS xdec64_3v512x8m81_0/RWL[16]
+ rcol4_512_3v512x8m81_0/WL[38] rcol4_512_3v512x8m81_0/WL[45] VSS xdec64_3v512x8m81_0/RWL[42]
+ VSS rcol4_512_3v512x8m81_0/WL[31] VSS VSS xdec64_3v512x8m81_0/RWL[27] xdec64_3v512x8m81_0/RWL[20]
+ rcol4_512_3v512x8m81_0/WL[58] rcol4_512_3v512x8m81_0/WL[60] rcol4_512_3v512x8m81_0/WL[62]
+ xdec64_3v512x8m81_0/RWL[29] xdec64_3v512x8m81_0/RWL[51] xdec64_3v512x8m81_0/RWL[55]
+ xdec64_3v512x8m81_0/RWL[57] VSS xdec64_3v512x8m81_0/RWL[7] rcol4_512_3v512x8m81_0/WL[8]
+ xdec64_3v512x8m81_0/RWL[5] VSS rcol4_512_3v512x8m81_0/WL[13] rcol4_512_3v512x8m81_0/WL[6]
+ rcol4_512_3v512x8m81_0/tblhl rcol4_512_3v512x8m81_0/GWE xdec64_3v512x8m81_0/RWL[11]
+ rcol4_512_3v512x8m81_0/din[7] rcol4_512_3v512x8m81_0/q[5] rcol4_512_3v512x8m81_0/q[6]
+ rcol4_512_3v512x8m81_0/q[7] rcol4_512_3v512x8m81_0/din[5] rcol4_512_3v512x8m81_0/din[6]
+ rcol4_512_3v512x8m81_0/q[4] rcol4_512_3v512x8m81_0/pcb[7] rcol4_512_3v512x8m81_0/pcb[4]
+ WEN[7] WEN[4] rcol4_512_3v512x8m81_0/pcb[5] WEN[6] WEN[5] D[7] control_3v512x8_3v512x8m81_0/RYS[1]
+ xdec64_3v512x8m81_0/RWL[21] xdec64_3v512x8m81_0/RWL[15] control_3v512x8_3v512x8m81_0/RYS[6]
+ xdec64_3v512x8m81_0/men xdec64_3v512x8m81_0/RWL[19] xdec64_3v512x8m81_0/RWL[8] xdec64_3v512x8m81_0/RWL[59]
+ VSS rcol4_512_3v512x8m81_0/saout_R_m2_3v512x8m81_1/sa_3v512x8m81_0/pcb xdec64_3v512x8m81_0/RWL[58]
+ Q[6] xdec64_3v512x8m81_0/RWL[6] xdec64_3v512x8m81_0/RWL[43] control_3v512x8_3v512x8m81_0/RYS[7]
+ xdec64_3v512x8m81_0/RWL[1] control_3v512x8_3v512x8m81_0/RYS[2] xdec64_3v512x8m81_0/RWL[36]
+ xdec64_3v512x8m81_0/RWL[22] xdec64_3v512x8m81_0/RWL[10] xdec64_3v512x8m81_0/RWL[61]
+ xdec64_3v512x8m81_0/RWL[46] xdec64_3v512x8m81_0/RWL[32] xdec64_3v512x8m81_0/RWL[60]
+ xdec64_3v512x8m81_0/RWL[9] control_3v512x8_3v512x8m81_0/RYS[0] xdec64_3v512x8m81_0/RWL[45]
+ xdec64_3v512x8m81_0/RWL[2] xdec64_3v512x8m81_0/RWL[39] xdec64_3v512x8m81_0/RWL[38]
+ xdec64_3v512x8m81_0/RWL[0] xdec64_3v512x8m81_0/RWL[24] xdec64_3v512x8m81_0/RWL[23]
+ xdec64_3v512x8m81_0/DRWL xdec64_3v512x8m81_0/RWL[12] D[5] control_3v512x8_3v512x8m81_0/IGWEN
+ rcol4_512_3v512x8m81_0/saout_R_m2_3v512x8m81_1/sa_3v512x8m81_0/pcb xdec64_3v512x8m81_0/RWL[48]
+ xdec64_3v512x8m81_0/RWL[62] control_3v512x8_3v512x8m81_0/RYS[4] xdec64_3v512x8m81_0/RWL[47]
+ xdec64_3v512x8m81_0/RWL[4] xdec64_3v512x8m81_0/RWL[26] xdec64_3v512x8m81_0/RWL[41]
+ Q[7] Q[4] xdec64_3v512x8m81_0/RWL[3] xdec64_3v512x8m81_0/RWL[40] xdec64_3v512x8m81_0/RWL[25]
+ control_3v512x8_3v512x8m81_0/RYS[3] Q[5] xdec64_3v512x8m81_0/RWL[14] control_3v512x8_3v512x8m81_0/RYS[5]
+ xdec64_3v512x8m81_0/RWL[49] xdec64_3v512x8m81_0/RWL[13] xdec64_3v512x8m81_0/RWL[18]
+ xdec64_3v512x8m81_0/RWL[34] xdec64_3v512x8m81_0/RWL[63] xdec64_3v512x8m81_0/RWL[17]
+ VSS VDD rcol4_512_3v512x8m81
Xxdec64_3v512x8m81_0 xdec64_3v512x8m81_0/DRWL xdec64_3v512x8m81_0/RWL[34] xdec64_3v512x8m81_0/RWL[35]
+ xdec64_3v512x8m81_0/RWL[36] xdec64_3v512x8m81_0/RWL[37] xdec64_3v512x8m81_0/RWL[38]
+ xdec64_3v512x8m81_0/RWL[39] xdec64_3v512x8m81_0/RWL[40] xdec64_3v512x8m81_0/RWL[42]
+ xdec64_3v512x8m81_0/RWL[44] xdec64_3v512x8m81_0/RWL[47] xdec64_3v512x8m81_0/RWL[49]
+ xdec64_3v512x8m81_0/RWL[50] xdec64_3v512x8m81_0/RWL[51] xdec64_3v512x8m81_0/RWL[52]
+ xdec64_3v512x8m81_0/RWL[53] xdec64_3v512x8m81_0/RWL[54] xdec64_3v512x8m81_0/RWL[55]
+ xdec64_3v512x8m81_0/RWL[56] xdec64_3v512x8m81_0/RWL[57] xdec64_3v512x8m81_0/RWL[58]
+ xdec64_3v512x8m81_0/RWL[60] xdec64_3v512x8m81_0/RWL[62] xdec64_3v512x8m81_0/LWL[62]
+ xdec64_3v512x8m81_0/LWL[61] xdec64_3v512x8m81_0/LWL[57] xdec64_3v512x8m81_0/LWL[55]
+ xdec64_3v512x8m81_0/LWL[53] xdec64_3v512x8m81_0/LWL[52] xdec64_3v512x8m81_0/LWL[50]
+ xdec64_3v512x8m81_0/LWL[49] xdec64_3v512x8m81_0/LWL[48] xdec64_3v512x8m81_0/LWL[37]
+ xdec64_3v512x8m81_0/LWL[35] xdec64_3v512x8m81_0/DLWL xdec64_3v512x8m81_0/LWL[19]
+ xdec64_3v512x8m81_0/LWL[20] xdec64_3v512x8m81_0/LWL[21] xdec64_3v512x8m81_0/LWL[22]
+ xdec64_3v512x8m81_0/LWL[26] xdec64_3v512x8m81_0/LWL[10] xdec64_3v512x8m81_0/LWL[12]
+ xdec64_3v512x8m81_0/LWL[14] xdec64_3v512x8m81_0/LWL[15] xdec64_3v512x8m81_0/LWL[17]
+ xdec64_3v512x8m81_0/LWL[18] xdec64_3v512x8m81_0/LWL[5] xdec64_3v512x8m81_0/LWL[4]
+ xdec64_3v512x8m81_0/LWL[3] xdec64_3v512x8m81_0/LWL[8] xdec64_3v512x8m81_0/LWL[9]
+ xdec64_3v512x8m81_0/LWL[6] xdec64_3v512x8m81_0/LWL[7] xdec64_3v512x8m81_0/RWL[31]
+ xdec64_3v512x8m81_0/RWL[25] xdec64_3v512x8m81_0/RWL[6] xdec64_3v512x8m81_0/RWL[4]
+ xdec64_3v512x8m81_0/RWL[5] xdec64_3v512x8m81_0/RWL[7] xdec64_3v512x8m81_0/RWL[8]
+ xdec64_3v512x8m81_0/RWL[10] xdec64_3v512x8m81_0/RWL[12] xdec64_3v512x8m81_0/RWL[13]
+ xdec64_3v512x8m81_0/RWL[14] xdec64_3v512x8m81_0/RWL[15] xdec64_3v512x8m81_0/xb[0]
+ xdec64_3v512x8m81_0/xb[1] xdec64_3v512x8m81_0/xb[2] xdec64_3v512x8m81_0/xb[3] xdec64_3v512x8m81_0/xa[7]
+ xdec64_3v512x8m81_0/xa[6] xdec64_3v512x8m81_0/xa[5] xdec64_3v512x8m81_0/xa[4] xdec64_3v512x8m81_0/xa[0]
+ xdec64_3v512x8m81_0/men xdec64_3v512x8m81_0/xa[3] xdec64_3v512x8m81_0/xa[2] xdec64_3v512x8m81_0/xa[1]
+ xdec64_3v512x8m81_0/xc[0] xdec64_3v512x8m81_0/xc[1] xdec64_3v512x8m81_0/LWL[24]
+ xdec64_3v512x8m81_0/RWL[59] xdec64_3v512x8m81_0/LWL[45] xdec64_3v512x8m81_0/LWL[29]
+ xdec64_3v512x8m81_0/LWL[63] xdec64_3v512x8m81_0/RWL[28] xdec64_3v512x8m81_0/RWL[23]
+ xdec64_3v512x8m81_0/LWL[46] xdec64_3v512x8m81_0/LWL[43] xdec64_3v512x8m81_0/RWL[26]
+ xdec64_3v512x8m81_0/LWL[27] xdec64_3v512x8m81_0/RWL[45] xdec64_3v512x8m81_0/LWL[44]
+ xdec64_3v512x8m81_0/RWL[24] lcol4_512_3v512x8m81_0/WL[59] xdec64_3v512x8m81_0/RWL[2]
+ xdec64_3v512x8m81_0/xdec32_468_3v512x8m81_0/LWL[30] xdec64_3v512x8m81_0/LWL[42]
+ xdec64_3v512x8m81_0/LWL[33] xdec64_3v512x8m81_0/RWL[3] xdec64_3v512x8m81_0/LWL[13]
+ xdec64_3v512x8m81_0/RWL[22] xdec64_3v512x8m81_0/RWL[11] xdec64_3v512x8m81_0/RWL[21]
+ xdec64_3v512x8m81_0/RWL[63] xdec64_3v512x8m81_0/LWL[32] xdec64_3v512x8m81_0/LWL[2]
+ xdec64_3v512x8m81_0/RWL[29] xdec64_3v512x8m81_0/RWL[0] xdec64_3v512x8m81_0/LWL[41]
+ xdec64_3v512x8m81_0/LWL[60] xdec64_3v512x8m81_0/LWL[40] xdec64_3v512x8m81_0/LWL[25]
+ xdec64_3v512x8m81_0/RWL[20] xdec64_3v512x8m81_0/LWL[1] xdec64_3v512x8m81_0/RWL[43]
+ xdec64_3v512x8m81_0/LWL[0] xdec64_3v512x8m81_0/RWL[32] xdec64_3v512x8m81_0/RWL[30]
+ xdec64_3v512x8m81_0/LWL[58] xdec64_3v512x8m81_0/LWL[38] xdec64_3v512x8m81_0/LWL[51]
+ xdec64_3v512x8m81_0/RWL[48] xdec64_3v512x8m81_0/RWL[18] VDD xdec64_3v512x8m81_0/LWL[59]
+ xdec64_3v512x8m81_0/LWL[30] xdec64_3v512x8m81_0/RWL[33] xdec64_3v512x8m81_0/RWL[1]
+ xdec64_3v512x8m81_0/LWL[56] xdec64_3v512x8m81_0/LWL[11] xdec64_3v512x8m81_0/LWL[36]
+ xdec64_3v512x8m81_0/RWL[19] xdec64_3v512x8m81_0/RWL[9] xdec64_3v512x8m81_0/RWL[61]
+ xdec64_3v512x8m81_0/RWL[46] xdec64_3v512x8m81_0/LWL[16] xdec64_3v512x8m81_0/RWL[17]
+ xdec64_3v512x8m81_0/RWL[27] xdec64_3v512x8m81_0/LWL[39] xdec64_3v512x8m81_0/LWL[28]
+ xdec64_3v512x8m81_0/LWL[47] xdec64_3v512x8m81_0/RWL[16] xdec64_3v512x8m81_0/LWL[23]
+ xdec64_3v512x8m81_0/LWL[54] xdec64_3v512x8m81_0/LWL[34] VSS xdec64_3v512x8m81_0/LWL[31]
+ xdec64_3v512x8m81_0/RWL[41] xdec64_3v512x8m81
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
X0 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 VDD I ZN VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7 VSS I ZN VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X9 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X13 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VNW VPW VSS
X0 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS I ZN VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD I ZN VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
X0 VDD a_572_375# a_484_472# VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt lvlshift_down VDD DVDD AH DVSS YL
Xgf180mcu_fd_sc_mcu7t5v0__inv_8_0 AH gf180mcu_fd_sc_mcu7t5v0__inv_8_0/ZN DVDD DVDD
+ DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xgf180mcu_fd_sc_mcu7t5v0__antenna_0 AH DVDD DVDD DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xgf180mcu_fd_sc_mcu7t5v0__inv_12_0 gf180mcu_fd_sc_mcu7t5v0__inv_8_0/ZN YL VDD VDD
+ DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__inv_12
Xgf180mcu_fd_sc_mcu7t5v0__fillcap_8_0 DVDD DVDD DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

.subckt pmos_6p0_GUW2N9 a_50_n324# w_n378_n586# a_n148_n324# a_n60_n368#
X0 a_50_n324# a_n60_n368# a_n148_n324# w_n378_n586# pfet_05v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.55u
.ends

.subckt nmos_6p0_BUMBUS a_n302_n300# a_n70_n168# a_n158_n76# a_70_n76#
X0 a_70_n76# a_n70_n168# a_n158_n76# a_n302_n300# nfet_05v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt pmos_6p0_MUW2NR a_n52_n524# w_n480_n786# a_162_n524# a_n162_n568# a_n250_n524#
+ a_52_n568#
X0 a_n52_n524# a_n162_n568# a_n250_n524# w_n480_n786# pfet_05v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.55u
X1 a_162_n524# a_52_n568# a_n52_n524# w_n480_n786# pfet_05v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.55u
.ends

.subckt nmos_6p0_BUMBJU a_n158_n276# a_n302_n500# a_n70_n368# a_70_n276#
X0 a_70_n276# a_n70_n368# a_n158_n276# a_n302_n500# nfet_05v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt std_inverter VDD Vin Vout VSS
XXM0 Vout VDD VDD Vin VDD Vin pmos_6p0_MUW2NR
XXM1 VSS VSS Vin Vout nmos_6p0_BUMBJU
.ends

.subckt std_buffer VDD Vin Vout VSS
XXM2 X0/Vin VDD VDD Vin pmos_6p0_GUW2N9
XXM3 VSS Vin VSS X0/Vin nmos_6p0_BUMBUS
XX0 VDD X0/Vin Vout VSS std_inverter
.ends

.subckt nmos_6p0_BJPB5U a_n70_n268# a_n158_n224# a_70_n224# a_n302_n400#
X0 a_70_n224# a_n70_n268# a_n158_n224# a_n302_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt pmos_6p0_EYEQQM a_n304_n268# a_n622_n176# a_234_n176# a_n408_n176# a_124_n268#
+ a_n732_n268# w_n1050_n486# a_n518_n268# a_n90_n268# a_662_n176# a_n820_n176# a_448_n176#
+ a_n194_n176# a_552_n268# a_20_n176# a_338_n268#
X0 a_448_n176# a_338_n268# a_234_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X1 a_n194_n176# a_n304_n268# a_n408_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X2 a_n408_n176# a_n518_n268# a_n622_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X3 a_662_n176# a_552_n268# a_448_n176# w_n1050_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.55u
X4 a_20_n176# a_n90_n268# a_n194_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X5 a_n622_n176# a_n732_n268# a_n820_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.55u
X6 a_234_n176# a_124_n268# a_20_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
.ends

.subckt nmos_6p0_B4TB5U a_n70_n268# a_70_n176# a_n158_n176# a_n302_n400#
X0 a_70_n176# a_n70_n268# a_n158_n176# a_n302_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt pmos_6p0_CYEQN4 a_n138_n176# a_60_n176# a_n50_n268# w_n368_n486#
X0 a_60_n176# a_n50_n268# a_n138_n176# w_n368_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.55u
.ends

.subckt nmos_6p0_BJXXPT a_662_n268# a_n314_n268# a_n70_n268# a_n418_n224# a_n1034_n400#
+ a_n174_n224# a_802_n224# a_n802_n268# a_n890_n224# a_n662_n224# a_418_n268# a_174_n268#
+ a_558_n224# a_314_n224# a_70_n224# a_n558_n268#
X0 a_n662_n224# a_n802_n268# a_n890_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X1 a_n174_n224# a_n314_n268# a_n418_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X2 a_802_n224# a_662_n268# a_558_n224# a_n1034_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X3 a_n418_n224# a_n558_n268# a_n662_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X4 a_70_n224# a_n70_n268# a_n174_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X5 a_314_n224# a_174_n268# a_70_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X6 a_558_n224# a_418_n268# a_314_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
.ends

.subckt ppolyf_u_1k_6p0_TRTT7C a_7600_n2622# a_5360_2500# a_2560_n2622# a_3120_n2622#
+ a_n5280_2500# a_8720_n2622# a_4800_2500# a_12080_n2622# a_3680_n2622# a_n8080_n2622#
+ a_600_2500# a_4240_n2622# a_n4720_2500# a_9840_n2622# a_6200_2500# a_5640_2500#
+ a_n1640_n2622# a_n10040_n2622# a_5360_n2622# a_n6120_2500# a_11800_n2622# a_880_2500#
+ a_n2200_n2622# a_n5560_2500# a_n240_2500# a_n7800_n2622# a_n240_n2622# a_n2760_n2622#
+ a_n11160_n2622# a_6480_n2622# a_7040_2500# a_6480_2500# a_n3320_n2622# a_7040_n2622#
+ a_n8920_n2622# a_n3880_n2622# a_n12280_n2622# a_5920_2500# a_n4440_n2622# a_8160_n2622#
+ a_n6400_2500# a_n5840_2500# a_n520_2500# a_n5000_n2622# a_1160_2500# a_7320_2500#
+ a_n5560_n2622# a_6760_2500# a_9280_n2622# a_320_n2622# a_n1080_2500# a_10120_n2622#
+ a_1720_n2622# a_n6120_n2622# a_n7240_2500# a_880_n2622# a_n1080_n2622# a_n6680_2500#
+ a_10680_n2622# a_n6680_n2622# a_8160_2500# a_11240_n2622# a_2840_n2622# a_n7240_n2622#
+ a_2000_2500# a_n800_2500# a_3400_n2622# a_1440_2500# a_n8080_2500# a_7600_2500#
+ a_n1360_2500# a_n8360_n2622# a_3960_n2622# a_4520_n2622# a_n7520_2500# a_n6960_2500#
+ a_2280_2500# a_n9480_n2622# a_n10040_2500# a_9000_2500# a_8440_2500# a_5640_n2622#
+ a_n1920_n2622# a_n10320_n2622# a_7880_2500# a_10120_2500# a_6200_n2622# a_1720_2500#
+ a_n8360_2500# a_n10880_n2622# a_n520_n2622# a_n2200_2500# a_1160_n2622# a_n1640_2500#
+ a_n11440_n2622# a_6760_n2622# a_9280_2500# a_n3600_n2622# a_n7800_2500# a_n12000_n2622#
+ a_7320_n2622# a_3120_2500# a_n10320_2500# a_2560_2500# a_2280_n2622# a_7880_n2622#
+ a_n3040_2500# a_8720_2500# a_n2480_2500# a_n4720_n2622# a_8440_n2622# a_10400_2500#
+ a_n9200_2500# a_n12492_n2834# a_n8640_2500# a_40_n2622# a_9000_n2622# a_n1920_2500#
+ a_n11160_2500# a_n5840_n2622# a_9560_n2622# a_9560_2500# a_10400_n2622# a_600_n2622#
+ a_11240_2500# a_n6400_n2622# a_3400_2500# a_10680_2500# a_n9480_2500# a_n10600_2500#
+ a_10960_n2622# a_2840_2500# a_n1360_n2622# a_5080_n2622# a_n3320_2500# a_n6960_n2622#
+ a_11520_n2622# a_n2760_2500# a_n7520_n2622# a_n8920_2500# a_12080_2500# a_n2480_n2622#
+ a_n12000_2500# a_4240_2500# a_3680_2500# a_n11440_2500# a_n3040_n2622# a_n10880_2500#
+ a_n4160_2500# a_n8640_n2622# a_9840_2500# a_11520_2500# a_4800_n2622# a_10960_2500#
+ a_n9200_n2622# a_n9760_2500# a_n4160_n2622# a_5080_2500# a_40_2500# a_n3600_2500#
+ a_n9760_n2622# a_n12280_2500# a_n10600_n2622# a_5920_n2622# a_n5280_n2622# a_4520_2500#
+ a_3960_2500# a_n5000_2500# a_n11720_2500# a_1440_n2622# a_320_2500# a_n800_n2622#
+ a_n4440_2500# a_n11720_n2622# a_n3880_2500# a_11800_2500# a_2000_n2622#
X0 a_n6400_2500# a_n6400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X1 a_n3320_2500# a_n3320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X2 a_1720_2500# a_1720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X3 a_7040_2500# a_7040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X4 a_n5840_2500# a_n5840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X5 a_9560_2500# a_9560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X6 a_n10040_2500# a_n10040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X7 a_5080_2500# a_5080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X8 a_n3880_2500# a_n3880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X9 a_n1360_2500# a_n1360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X10 a_2000_2500# a_2000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X11 a_4520_2500# a_4520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X12 a_n10600_2500# a_n10600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X13 a_n9200_2500# a_n9200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X14 a_n6120_2500# a_n6120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X15 a_11520_2500# a_11520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X16 a_12080_2500# a_12080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X17 a_n8640_2500# a_n8640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X18 a_n4160_2500# a_n4160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X19 a_2560_2500# a_2560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X20 a_n6680_2500# a_n6680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X21 a_7320_2500# a_7320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X22 a_9840_2500# a_9840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X23 a_n10320_2500# a_n10320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X24 a_n2200_2500# a_n2200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X25 a_5360_2500# a_5360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X26 a_n1640_2500# a_n1640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X27 a_4800_2500# a_4800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X28 a_7880_2500# a_7880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X29 a_n10880_2500# a_n10880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X30 a_n9480_2500# a_n9480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X31 a_n8920_2500# a_n8920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X32 a_11800_2500# a_11800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X33 a_2840_2500# a_2840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X34 a_n4440_2500# a_n4440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X35 a_8160_2500# a_8160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X36 a_n11160_2500# a_n11160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X37 a_n6960_2500# a_n6960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X38 a_320_2500# a_320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X39 a_7600_2500# a_7600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X40 a_n5000_2500# a_n5000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X41 a_n2480_2500# a_n2480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X42 a_n1920_2500# a_n1920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X43 a_3120_2500# a_3120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X44 a_5640_2500# a_5640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X45 a_n9760_2500# a_n9760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X46 a_n7240_2500# a_n7240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X47 a_880_2500# a_880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X48 a_10120_2500# a_10120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X49 a_1160_2500# a_1160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X50 a_3680_2500# a_3680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X51 a_n5280_2500# a_n5280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X52 a_n240_2500# a_n240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X53 a_40_2500# a_40_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X54 a_n7800_2500# a_n7800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X55 a_n4720_2500# a_n4720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X56 a_8440_2500# a_8440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X57 a_10680_2500# a_10680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X58 a_n11440_2500# a_n11440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X59 a_600_2500# a_600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X60 a_n2760_2500# a_n2760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X61 a_n800_2500# a_n800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X62 a_3400_2500# a_3400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X63 a_6480_2500# a_6480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X64 a_n8080_2500# a_n8080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X65 a_5920_2500# a_5920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X66 a_n12000_2500# a_n12000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X67 a_n7520_2500# a_n7520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X68 a_10400_2500# a_10400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X69 a_1440_2500# a_1440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X70 a_3960_2500# a_3960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X71 a_n5560_2500# a_n5560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X72 a_n3040_2500# a_n3040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X73 a_n520_2500# a_n520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X74 a_6200_2500# a_6200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X75 a_9280_2500# a_9280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X76 a_10960_2500# a_10960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X77 a_n12280_2500# a_n12280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X78 a_8720_2500# a_8720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X79 a_n11720_2500# a_n11720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X80 a_n3600_2500# a_n3600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X81 a_n1080_2500# a_n1080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X82 a_4240_2500# a_4240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X83 a_6760_2500# a_6760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X84 a_n8360_2500# a_n8360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X85 a_9000_2500# a_9000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X86 a_11240_2500# a_11240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X87 a_2280_2500# a_2280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
.ends

.subckt pmos_6p0_HUEQQM a_375_n176# a_265_n268# a_n810_n268# a_n596_n268# a_803_n176#
+ a_n272_n176# a_589_n176# a_161_n176# a_693_n268# a_n58_n176# a_479_n268# a_51_n268#
+ a_n382_n268# w_n1128_n486# a_n168_n268# a_n898_n176# a_n700_n176# a_n486_n176#
X0 a_375_n176# a_265_n268# a_161_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X1 a_n272_n176# a_n382_n268# a_n486_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X2 a_n700_n176# a_n810_n268# a_n898_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.55u
X3 a_589_n176# a_479_n268# a_375_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X4 a_n486_n176# a_n596_n268# a_n700_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X5 a_161_n176# a_51_n268# a_n58_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.545p ps=2.545u w=2u l=0.55u
X6 a_n58_n176# a_n168_n268# a_n272_n176# w_n1128_n486# pfet_05v0 ad=0.545p pd=2.545u as=0.52p ps=2.52u w=2u l=0.55u
X7 a_803_n176# a_693_n268# a_589_n176# w_n1128_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.55u
.ends

.subckt reduction_mirror VDD Vout VSS
Xnmos_6p0_BJPB5U_0 m2_1393_n86# VSS m2_3858_n195# VSS nmos_6p0_BJPB5U
Xpmos_6p0_EYEQQM_0 m2_4433_1027# VDD VDD m2_4433_1027# m2_4433_1027# m2_4433_1027#
+ VDD m2_4433_1027# m2_4433_1027# VDD m2_4433_1027# m2_4433_1027# VDD m2_4433_1027#
+ m2_4433_1027# m2_4433_1027# pmos_6p0_EYEQQM
XXM0 m1_2517_n836# VSS m2_607_119# VSS nmos_6p0_B4TB5U
XXM1 m2_3432_1017# m2_1393_n86# m2_607_119# VDD pmos_6p0_CYEQN4
Xpmos_6p0_CYEQN4_0 m2_6726_1023# Vout m2_3858_n195# VDD pmos_6p0_CYEQN4
XXM3 m2_607_119# m2_921_1004# m2_607_119# VDD pmos_6p0_CYEQN4
XXM4 VDD m2_3432_1017# m2_921_1004# VDD pmos_6p0_CYEQN4
XXM7 VDD m2_6726_1023# m2_4433_1027# VDD pmos_6p0_CYEQN4
XXM9 m2_3858_n195# m2_4433_1027# m2_3858_n195# VDD pmos_6p0_CYEQN4
Xnmos_6p0_BJXXPT_0 m2_1393_n86# m2_1393_n86# m2_1393_n86# m2_1393_n86# VSS VSS VSS
+ m2_1393_n86# m2_1393_n86# VSS m2_1393_n86# m2_1393_n86# m2_1393_n86# VSS m2_1393_n86#
+ m2_1393_n86# nmos_6p0_BJXXPT
Xppolyf_u_1k_6p0_TRTT7C_0 m1_20155_n6001# m1_18197_n836# m1_15115_n6001# m1_15675_n6001#
+ m1_7557_n836# m1_21275_n6001# m1_17637_n836# m1_24635_n6001# m1_16235_n6001# m1_4475_n6001#
+ m1_13157_n836# m1_16795_n6001# m1_8117_n836# m1_22395_n6001# m1_18757_n836# m1_18197_n836#
+ m1_11195_n6001# m1_2795_n6001# m1_17915_n6001# m1_6437_n836# m1_24635_n6001# m1_13717_n836#
+ m1_10635_n6001# m1_6997_n836# m1_12597_n836# m1_5035_n6001# m1_12315_n6001# m1_10075_n6001#
+ m1_1675_n6001# m1_19035_n6001# m1_19877_n836# m1_19317_n836# m1_9515_n6001# m1_19595_n6001#
+ m1_3915_n6001# m1_8955_n6001# m1_555_n6001# m1_18757_n836# m1_8395_n6001# m1_20715_n6001#
+ m1_6437_n836# m1_6997_n836# m1_12037_n836# m1_7835_n6001# m1_13717_n836# m1_19877_n836#
+ m1_7275_n6001# m1_19317_n836# m1_21835_n6001# m1_12875_n6001# m1_11477_n836# m1_22955_n6001#
+ m1_14555_n6001# m1_6715_n6001# m1_5317_n836# m1_13435_n6001# m1_11755_n6001# m1_5877_n836#
+ m1_23515_n6001# m1_6155_n6001# m1_20997_n836# m1_24075_n6001# m1_15675_n6001# m1_5595_n6001#
+ m1_14837_n836# m1_12037_n836# m1_16235_n6001# m1_14277_n836# m1_4757_n836# m1_20437_n836#
+ m1_11477_n836# m1_4475_n6001# m1_16795_n6001# m1_17355_n6001# m1_5317_n836# m1_5877_n836#
+ m1_14837_n836# m1_3355_n6001# m1_2517_n836# m1_21557_n836# m1_20997_n836# m1_18475_n6001#
+ m1_10635_n6001# m1_2235_n6001# m1_20437_n836# m1_22677_n836# m1_19035_n6001# m1_14277_n836#
+ m1_4197_n836# m1_1675_n6001# m1_12315_n6001# m1_10357_n836# m1_13995_n6001# m1_10917_n836#
+ m1_1115_n6001# m1_19595_n6001# m1_22117_n836# m1_8955_n6001# m1_4757_n836# m1_555_n6001#
+ m1_20155_n6001# m1_15957_n836# m1_2517_n836# m1_15397_n836# m1_15115_n6001# m1_20715_n6001#
+ m1_9797_n836# m1_21557_n836# m1_10357_n836# m1_7835_n6001# m1_21275_n6001# m1_23237_n836#
+ m1_3637_n836# VSS m1_4197_n836# m1_12875_n6001# m1_21835_n6001# m1_10917_n836# m1_1397_n836#
+ m1_6715_n6001# m1_22395_n6001# m1_22117_n836# m1_22955_n6001# m1_13435_n6001# m1_23797_n836#
+ m1_6155_n6001# m1_15957_n836# m1_23237_n836# m1_3077_n836# m1_1957_n836# m1_23515_n6001#
+ m1_15397_n836# m1_11195_n6001# m1_17915_n6001# m1_9237_n836# m1_5595_n6001# m1_24075_n6001#
+ m1_9797_n836# m1_5035_n6001# m1_3637_n836# VDD m1_10075_n6001# m1_837_n836# m1_17077_n836#
+ m1_16517_n836# m1_1397_n836# m1_9515_n6001# m1_1957_n836# m1_8677_n836# m1_3915_n6001#
+ m1_22677_n836# m1_24357_n836# m1_17355_n6001# m1_23797_n836# m1_3355_n6001# m1_3077_n836#
+ m1_8395_n6001# m1_17637_n836# m1_12597_n836# m1_9237_n836# m1_2795_n6001# VSS m1_2235_n6001#
+ m1_18475_n6001# m1_7275_n6001# m1_17077_n836# m1_16517_n836# m1_7557_n836# m1_837_n836#
+ m1_13995_n6001# m1_13157_n836# m1_11755_n6001# m1_8117_n836# m1_1115_n6001# m1_8677_n836#
+ m1_24357_n836# m1_14555_n6001# ppolyf_u_1k_6p0_TRTT7C
Xpmos_6p0_HUEQQM_0 m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004#
+ VDD VDD VDD m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# VDD
+ m2_921_1004# m2_921_1004# VDD m2_921_1004# pmos_6p0_HUEQQM
.ends

.subckt mim_2p0fF_8KW78G m4_n1220_n1120# m4_n1100_n1000#
X0 m4_n1100_n1000# m4_n1220_n1120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=10u
.ends

.subckt large_mimcap In VSS
XXC1[0|0] VSS In mim_2p0fF_8KW78G
XXC1[1|0] VSS In mim_2p0fF_8KW78G
XXC1[2|0] VSS In mim_2p0fF_8KW78G
XXC1[0|1] VSS In mim_2p0fF_8KW78G
XXC1[1|1] VSS In mim_2p0fF_8KW78G
XXC1[2|1] VSS In mim_2p0fF_8KW78G
XXC1[0|2] VSS In mim_2p0fF_8KW78G
XXC1[1|2] VSS In mim_2p0fF_8KW78G
XXC1[2|2] VSS In mim_2p0fF_8KW78G
.ends

.subckt pmos_6p0_UXEQNM a_n60_n168# a_n148_n76# w_n378_n386# a_50_n76#
X0 a_50_n76# a_n60_n168# a_n148_n76# w_n378_n386# pfet_05v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt nmos_6p0_L3YBEV a_n188_n724# a_100_n724# a_n332_n900# a_n100_n768#
X0 a_100_n724# a_n100_n768# a_n188_n724# a_n332_n900# nfet_05v0 ad=3.08p pd=14.88u as=3.08p ps=14.88u w=7u l=1u
.ends

.subckt pmos_6p0_9YEQN4 a_50_n576# w_n378_n886# a_n148_n576# a_n60_n668#
X0 a_50_n576# a_n60_n668# a_n148_n576# w_n378_n886# pfet_05v0 ad=2.64p pd=12.88u as=2.64p ps=12.88u w=6u l=0.55u
.ends

.subckt pmos_6p0_9859UL a_n288_n26# a_n200_n118# a_200_n26# w_n518_n336#
X0 a_200_n26# a_n200_n118# a_n288_n26# w_n518_n336# pfet_05v0 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=2u
.ends

.subckt schmitt_inverter VDD VSS Vin Vout
Xpmos_6p0_UXEQNM_0 Vin m1_1072_n872# VDD Vout pmos_6p0_UXEQNM
XX6 m1_1243_n1927# VDD VSS Vout nmos_6p0_L3YBEV
Xnmos_6p0_BJPB5U_0 Vin m1_1243_n1927# Vout VSS nmos_6p0_BJPB5U
XXM1 m1_1072_n872# VDD VDD Vin pmos_6p0_9YEQN4
XXM3 Vin VSS m1_1243_n1927# VSS nmos_6p0_BJPB5U
XXM5 m1_1072_n872# Vout VSS VDD pmos_6p0_9859UL
.ends

.subckt simple_por VDD porb por VSS
Xstd_buffer_0 VDD X3/Vin por VSS std_buffer
XX0 VDD X1/In VSS reduction_mirror
XX1 X1/In VSS large_mimcap
XX2 VDD VSS X1/In X3/Vin schmitt_inverter
XX3 VDD X3/Vin porb VSS std_inverter
.ends

.subckt x018SRAM_cell1_dummy_3v256x8m81 m3_82_330# a_248_342# a_248_592# w_82_512#
+ a_62_178# m2_346_89# m2_134_89# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_82_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_82_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt new_dummyrow_unit_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89# 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
X018SRAM_cell1_dummy_3v256x8m81_10 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt new_dummyrowunit01_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
X018SRAM_cell1_dummy_3v256x8m81_10 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt x018SRAM_cell1_3v256x8m81 m3_82_330# a_248_342# a_248_592# a_62_178# w_30_512#
+ a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt x018SRAM_cell1_cutPC_3v256x8m81 m3_82_330# a_248_342# a_248_592# a_62_178#
+ w_30_512# a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt array16_256_dummy_01_3v256x8m81 018SRAM_cell1_cutPC_3v256x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_61/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_62/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_14/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_10/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_62/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_57/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_15/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_48/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_11/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_54/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_50/a_62_178#
+ VSS VDD 018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_31/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_12/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_59/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_2/a_62_178#
+ VSUBS
X018SRAM_cell1_cutPC_3v256x8m81_4 018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_5 018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_5/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_6 018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_8 018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_7 018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_7/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_9 018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_60 018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_50 018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_50/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_61 018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_61/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_51 018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_62 018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v256x8m81_62/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_62/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_52 018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_53 018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_53/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_31 018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_31/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_63 018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_10 018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_10/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_54 018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_54/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_11 018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_11/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_55 018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_12 018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_12/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_56 018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_13 018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_57 018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_57/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_14 018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_14/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_58 018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_48 018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_48/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_15 018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_15/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_59 018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_59/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_49 018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_49/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_0 018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v256x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_2 018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330# VSS
+ 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_2/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_3 018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_3/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
.ends

.subckt ldummy_3v256x4_3v256x8m81 array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
Xnew_dummyrow_unit_3v256x8m81_0 new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ VSUBS new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ new_dummyrow_unit_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_10 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_21 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_22 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_23 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_24 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_25 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_26 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_16 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_27 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_17 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_28 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_18 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_29 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_19 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xnew_dummyrowunit01_3v256x8m81_0 new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# new_dummyrowunit01_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_0 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD VSUBS
+ array16_256_dummy_01_3v256x8m81_0/VDD 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD VSUBS
+ array16_256_dummy_01_3v256x8m81_0/VDD 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xarray16_256_dummy_01_3v256x8m81_0 VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# VSUBS
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592#
+ VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342#
+ VSUBS VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512#
+ VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342#
+ VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# VSUBS
+ VSUBS VSUBS VSUBS array16_256_dummy_01_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_30 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_31 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_20 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt pmos_5p04310591302030_3v256x8m81 a_871_n45# D a_n252_n45# a_550_n45# a_229_n45#
+ w_n426_n86# a_390_n45# S a_n92_n45# a_1032_n45# a_1192_n45# a_711_n45# a_69_n45#
X0 D a_390_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X1 D a_n252_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.5566p ps=3.41u w=1.265u l=0.28u
X2 D a_69_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X3 S a_229_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X4 S a_550_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X5 S a_1192_n45# D w_n426_n86# pfet_03v3 ad=0.5566p pd=3.41u as=0.3289p ps=1.785u w=1.265u l=0.28u
X6 D a_1032_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X7 S a_n92_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X8 S a_871_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X9 D a_711_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
.ends

.subckt pmos_1p2$$45095980_3v256x8m81 a_697_n34# pmos_5p04310591302030_3v256x8m81_0/D
+ a_n106_n34# a_n266_n34# a_376_n34# a_1018_n34# a_1178_n34# a_55_n34# a_857_n34#
+ pmos_5p04310591302030_3v256x8m81_0/S a_536_n34# w_987_n66# a_215_n34#
Xpmos_5p04310591302030_3v256x8m81_0 a_857_n34# pmos_5p04310591302030_3v256x8m81_0/D
+ a_n266_n34# a_536_n34# a_215_n34# w_987_n66# a_376_n34# pmos_5p04310591302030_3v256x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34# a_55_n34# pmos_5p04310591302030_3v256x8m81
.ends

.subckt pmos_5p04310591302027_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302029_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.54067p pd=3.32u as=0.3159p ps=1.735u w=1.215u l=0.28u
.ends

.subckt nmos_1p2$$45100076_3v256x8m81 nmos_5p04310591302029_3v256x8m81_0/S nmos_5p04310591302029_3v256x8m81_0/D
+ a_118_n34# a_n41_n34# VSUBS
Xnmos_5p04310591302029_3v256x8m81_0 nmos_5p04310591302029_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302029_3v256x8m81_0/S VSUBS nmos_5p04310591302029_3v256x8m81
.ends

.subckt pmos_5p04310591302024_3v256x8m81 w_n286_n86# a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S
X0 D a_n112_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_369_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_209_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 D a_530_n44# S w_n286_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X4 S a_48_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46282796_3v256x8m81 pmos_5p04310591302024_3v256x8m81_0/S a_n126_n34#
+ a_195_n34# pmos_5p04310591302024_3v256x8m81_0/D a_516_n34# w_163_n66# a_355_n34#
+ a_34_n34#
Xpmos_5p04310591302024_3v256x8m81_0 w_163_n66# a_516_n34# pmos_5p04310591302024_3v256x8m81_0/D
+ a_n126_n34# a_195_n34# a_355_n34# a_34_n34# pmos_5p04310591302024_3v256x8m81_0/S
+ pmos_5p04310591302024_3v256x8m81
.ends

.subckt nmos_5p04310591302032_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.23585p pd=1.95u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_5p04310591302022_3v256x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.8382p ps=4.69u w=1.905u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=0.8382p pd=4.69u as=0.4953p ps=2.425u w=1.905u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
.ends

.subckt pmos_1p2$$46283820_3v256x8m81 a_536_n34# a_215_n34# a_697_n34# a_n106_n34#
+ a_n266_n34# pmos_5p04310591302022_3v256x8m81_0/S a_376_n34# w_984_n66# a_1018_n34#
+ a_1178_n34# a_55_n34# a_857_n34# pmos_5p04310591302022_3v256x8m81_0/D
Xpmos_5p04310591302022_3v256x8m81_0 pmos_5p04310591302022_3v256x8m81_0/D a_n266_n34#
+ a_536_n34# a_215_n34# w_984_n66# a_376_n34# pmos_5p04310591302022_3v256x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34# a_55_n34# a_857_n34# pmos_5p04310591302022_3v256x8m81
.ends

.subckt nmos_5p04310591302036_3v256x8m81 a_530_n44# D a_n112_n44# a_209_n44# a_369_n44#
+ a_48_n44# S VSUBS
X0 D a_n112_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_369_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.13913p ps=1.055u w=0.53u l=0.28u
X3 D a_530_n44# S VSUBS nfet_03v3 ad=0.2332p pd=1.94u as=0.13913p ps=1.055u w=0.53u l=0.28u
X4 S a_48_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt nmos_1p2$$45101100_3v256x8m81 a_195_n34# nmos_5p04310591302036_3v256x8m81_0/S
+ a_35_n34# a_516_n34# nmos_5p04310591302036_3v256x8m81_0/D a_n125_n34# a_356_n34#
+ VSUBS
Xnmos_5p04310591302036_3v256x8m81_0 a_516_n34# nmos_5p04310591302036_3v256x8m81_0/D
+ a_n125_n34# a_195_n34# a_356_n34# a_35_n34# nmos_5p04310591302036_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302036_3v256x8m81
.ends

.subckt nmos_5p04310591302033_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.28u
.ends

.subckt pmos_5p04310591302031_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4134p pd=2.11u as=0.6996p ps=4.06u w=1.59u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6996p pd=4.06u as=0.4134p ps=2.11u w=1.59u l=0.28u
.ends

.subckt pmos_1p2$$46287916_3v256x8m81 w_n133_n66# pmos_5p04310591302031_3v256x8m81_0/S
+ a_n42_n34# pmos_5p04310591302031_3v256x8m81_0/D a_118_n34#
Xpmos_5p04310591302031_3v256x8m81_0 pmos_5p04310591302031_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302031_3v256x8m81_0/S pmos_5p04310591302031_3v256x8m81
.ends

.subckt nmos_5p04310591302026_3v256x8m81 a_154_n44# D a_n168_n44# a_476_n44# a_798_n44#
+ a_314_n44# a_n8_n44# S a_636_n44# VSUBS
X0 S a_636_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_314_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_n168_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X3 S a_n8_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_798_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X5 D a_476_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X6 D a_154_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$45102124_3v256x8m81 a_140_n34# nmos_5p04310591302026_3v256x8m81_0/S
+ a_462_n34# a_n181_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v256x8m81_0/D
+ a_622_n34# a_n22_n34# VSUBS
Xnmos_5p04310591302026_3v256x8m81_0 a_140_n34# nmos_5p04310591302026_3v256x8m81_0/D
+ a_n181_n34# a_462_n34# a_784_n34# a_300_n34# a_n22_n34# nmos_5p04310591302026_3v256x8m81_0/S
+ a_622_n34# VSUBS nmos_5p04310591302026_3v256x8m81
.ends

.subckt pmos_5p04310591302035_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$46284844_3v256x8m81 w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S
+ pmos_5p04310591302035_3v256x8m81_0/D a_118_n34# a_n42_n34#
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S pmos_5p04310591302035_3v256x8m81
.ends

.subckt pmos_5p04310591302013_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46286892_3v256x8m81 w_n133_n66# pmos_5p04310591302013_3v256x8m81_0/D
+ a_251_n34# a_n70_n34# a_90_n34# pmos_5p04310591302013_3v256x8m81_0/S
Xpmos_5p04310591302013_3v256x8m81_0 pmos_5p04310591302013_3v256x8m81_0/D a_251_n34#
+ pmos_5p04310591302013_3v256x8m81_0/S a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302013_3v256x8m81
.ends

.subckt nmos_5p04310591302028_3v256x8m81 D a_64_n44# a_226_n44# a_386_n44# a_548_n44#
+ S a_n96_n44# VSUBS
X0 D a_548_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X1 S a_386_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_226_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X3 D a_n96_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X4 S a_64_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302025_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n85#
X0 D a_265_n44# S w_n230_n85# pfet_03v3 ad=0.9306p pd=5.11u as=0.55518p ps=2.64u w=2.115u l=0.28u
X1 D a_n56_n44# S w_n230_n85# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X2 S a_104_n44# D w_n230_n85# pfet_03v3 ad=0.55518p pd=2.64u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$46281772_3v256x8m81 pmos_5p04310591302025_3v256x8m81_0/S a_251_n34#
+ w_n133_n66# a_n70_n34# pmos_5p04310591302025_3v256x8m81_0/D a_90_n34#
Xpmos_5p04310591302025_3v256x8m81_0 pmos_5p04310591302025_3v256x8m81_0/D a_251_n34#
+ pmos_5p04310591302025_3v256x8m81_0/S a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302025_3v256x8m81
.ends

.subckt nmos_5p04310591302023_3v256x8m81 D a_n32_n44# a_136_n44# S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=92.8f pd=0.92u as=0.1576p ps=1.64u w=0.28u l=0.28u
X1 S a_136_n44# D VSUBS nfet_03v3 ad=0.159p pd=1.65u as=92.8f ps=0.92u w=0.28u l=0.28u
.ends

.subckt pmos_5p04310591302014_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46285868_3v256x8m81 w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S
+ pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_5p04310591302038_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.2464p pd=2u as=0.2464p ps=2u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302037_3v256x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X1 S a_662_n44# D VSUBS nfet_03v3 ad=0.5852p pd=3.54u as=0.3458p ps=1.85u w=1.33u l=0.28u
X2 D a_502_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X3 S a_20_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X4 D a_181_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X5 D a_n140_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.5852p ps=3.54u w=1.33u l=0.28u
.ends

.subckt nmos_1p2$$45103148_3v256x8m81 a_327_n34# a_n153_n34# a_488_n34# nmos_5p04310591302037_3v256x8m81_0/S
+ a_167_n34# a_6_n34# nmos_5p04310591302037_3v256x8m81_0/D a_648_n34# VSUBS
Xnmos_5p04310591302037_3v256x8m81_0 a_6_n34# nmos_5p04310591302037_3v256x8m81_0/D
+ a_167_n34# a_488_n34# a_648_n34# a_n153_n34# nmos_5p04310591302037_3v256x8m81_0/S
+ a_327_n34# VSUBS nmos_5p04310591302037_3v256x8m81
.ends

.subckt nmos_5p04310591302012_3v256x8m81 a_n83_n44# D a_77_n44# S a_237_n44# a_397_n44#
+ VSUBS
X0 S a_77_n44# D VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_397_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_237_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X3 D a_n83_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt sacntl_2_3v256x8m81 pcb se men pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81_2/S
+ vss vdd
Xpmos_1p2$$45095980_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S se nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S
+ vdd nmos_5p04310591302028_3v256x8m81_1/S vdd nmos_5p04310591302028_3v256x8m81_1/S
+ pmos_1p2$$45095980_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_0 vdd pmos_5p04310591302027_3v256x8m81_2/S pmos_5p04310591302027_3v256x8m81_0/S
+ vdd pmos_5p04310591302027_3v256x8m81_0/S pmos_5p04310591302027_3v256x8m81
Xnmos_1p2$$45100076_3v256x8m81_0 vss pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ vss nmos_1p2$$45100076_3v256x8m81
Xpmos_1p2$$46282796_3v256x8m81_0 vdd men men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ men vdd men men pmos_1p2$$46282796_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_1 vdd pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vss vdd pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_2 vdd pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81_2/S
+ vdd pmos_5p04310591302027_3v256x8m81_2/S pmos_5p04310591302027_3v256x8m81
Xnmos_5p04310591302032_3v256x8m81_0 nmos_5p04310591302032_3v256x8m81_0/D pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D vss vss nmos_5p04310591302032_3v256x8m81
Xpmos_1p2$$46283820_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pcb pmos_1p2$$46283820_3v256x8m81
Xnmos_1p2$$45101100_3v256x8m81_0 men vss men men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ men men vss nmos_1p2$$45101100_3v256x8m81
Xnmos_5p04310591302033_3v256x8m81_0 vss pmos_5p04310591302027_3v256x8m81_0/S pmos_5p04310591302038_3v256x8m81_0/S
+ vss nmos_5p04310591302033_3v256x8m81
Xpmos_1p2$$46287916_3v256x8m81_0 vdd vdd pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ nmos_5p04310591302032_3v256x8m81_0/D pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_1p2$$46287916_3v256x8m81
Xnmos_1p2$$45102124_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vss pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pcb pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vss nmos_1p2$$45102124_3v256x8m81
Xpmos_1p2$$46284844_3v256x8m81_0 vdd vdd pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81_1/S pmos_1p2$$46284844_3v256x8m81
Xpmos_1p2$$46286892_3v256x8m81_0 vdd nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302032_3v256x8m81_0/D
+ nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D vdd pmos_1p2$$46286892_3v256x8m81
Xnmos_5p04310591302028_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/D nmos_5p04310591302032_3v256x8m81_0/D
+ nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D
+ vss nmos_5p04310591302032_3v256x8m81_0/D vss nmos_5p04310591302028_3v256x8m81
Xpmos_1p2$$46281772_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S vdd pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ vdd pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_0 vss pmos_5p04310591302027_3v256x8m81_2/S pmos_5p04310591302027_3v256x8m81_0/S
+ pmos_5p04310591302027_3v256x8m81_0/S vss nmos_5p04310591302023_3v256x8m81
Xnmos_5p04310591302028_3v256x8m81_1 nmos_5p04310591302028_3v256x8m81_1/D pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D nmos_5p04310591302028_3v256x8m81_1/S
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D vss nmos_5p04310591302028_3v256x8m81
Xpmos_1p2$$46281772_3v256x8m81_1 pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ nmos_5p04310591302028_3v256x8m81_1/S vdd pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vdd pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_1p2$$46281772_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_1 vss pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vss pmos_5p04310591302027_3v256x8m81_1/S vss nmos_5p04310591302023_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_2 vss pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81_2/S
+ pmos_5p04310591302027_3v256x8m81_2/S vss nmos_5p04310591302023_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 vdd nmos_5p04310591302028_3v256x8m81_1/S vdd pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46285868_3v256x8m81
Xpmos_5p04310591302038_3v256x8m81_0 vdd pmos_5p04310591302027_3v256x8m81_0/S vdd pmos_5p04310591302038_3v256x8m81_0/S
+ pmos_5p04310591302038_3v256x8m81
Xnmos_1p2$$45103148_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D vss nmos_5p04310591302028_3v256x8m81_1/S
+ pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D vss nmos_1p2$$45103148_3v256x8m81
Xnmos_5p04310591302012_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S se nmos_5p04310591302028_3v256x8m81_1/S
+ vss nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S vss
+ nmos_5p04310591302012_3v256x8m81
X0 pmos_1p2$$46284844_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302027_3v256x8m81_1/S vss vss nfet_03v3 ad=0.2948p pd=2.22u as=0.2948p ps=2.22u w=0.67u l=0.28u
.ends

.subckt nmos_5p04310591302050_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# VSUBS
X0 D a_265_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S a_104_n44# D VSUBS nfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302044_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.451p pd=2.93u as=0.451p ps=2.93u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302047_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.8206p pd=4.61u as=0.8206p ps=4.61u w=1.865u l=0.28u
.ends

.subckt nmos_5p04310591302045_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt pmos_5p04310591302048_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.924p pd=5.08u as=0.924p ps=5.08u w=2.1u l=0.28u
.ends

.subckt nmos_5p04310591302046_3v256x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X1 S a_662_n44# D VSUBS nfet_03v3 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.28u
X2 D a_502_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X3 S a_20_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X4 D a_181_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X5 D a_n140_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.28u
.ends

.subckt pmos_5p04310591302049_3v256x8m81 a_20_n44# D a_181_n44# a_n140_n44# S a_341_n44#
+ a_503_n44# a_663_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.4664p pd=2.29u as=0.4576p ps=2.28u w=1.76u l=0.28u
X1 S a_20_n44# D w_n314_n86# pfet_03v3 ad=0.462p pd=2.285u as=0.4576p ps=2.28u w=1.76u l=0.28u
X2 D a_181_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.462p ps=2.285u w=1.76u l=0.28u
X3 D a_n140_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.7744p ps=4.4u w=1.76u l=0.28u
X4 S a_663_n44# D w_n314_n86# pfet_03v3 ad=0.7832p pd=4.41u as=0.4576p ps=2.28u w=1.76u l=0.28u
X5 D a_503_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.4664p ps=2.29u w=1.76u l=0.28u
.ends

.subckt pmos_5p04310591302051_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6877p pd=3.165u as=1.1638p ps=6.17u w=2.645u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1638p pd=6.17u as=0.6877p ps=3.165u w=2.645u l=0.28u
.ends

.subckt pmos_5p0431059130203_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_1p2$$171625516_3v256x8m81 a_n42_n34# pmos_5p0431059130203_3v256x8m81_0/S
+ pmos_5p0431059130203_3v256x8m81_0/w_n202_n86# a_118_n34# pmos_5p0431059130203_3v256x8m81_0/D
Xpmos_5p0431059130203_3v256x8m81_0 pmos_5p0431059130203_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# pmos_5p0431059130203_3v256x8m81_0/w_n202_n86# pmos_5p0431059130203_3v256x8m81_0/S
+ pmos_5p0431059130203_3v256x8m81
.ends

.subckt outbuf_oe_3v256x8m81 qp qn se q GWE vss vdd
Xnmos_5p04310591302050_3v256x8m81_0 pmos_5p04310591302013_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_0/D
+ vss nmos_5p04310591302050_3v256x8m81
Xnmos_5p04310591302044_3v256x8m81_0 vss pmos_5p04310591302047_3v256x8m81_0/S pmos_5p04310591302048_3v256x8m81_0/S
+ vss nmos_5p04310591302044_3v256x8m81
Xpmos_5p04310591302047_3v256x8m81_0 vdd GWE vdd pmos_5p04310591302047_3v256x8m81_0/S
+ pmos_5p04310591302047_3v256x8m81
Xnmos_5p04310591302033_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ vss vss nmos_5p04310591302033_3v256x8m81
Xnmos_5p04310591302045_3v256x8m81_0 vss pmos_5p04310591302047_3v256x8m81_0/S pmos_5p04310591302047_3v256x8m81_0/S
+ nmos_5p04310591302045_3v256x8m81_1/S vss nmos_5p04310591302045_3v256x8m81
Xnmos_5p04310591302045_3v256x8m81_1 pmos_5p04310591302051_3v256x8m81_0/D qn qn nmos_5p04310591302045_3v256x8m81_1/S
+ vss nmos_5p04310591302045_3v256x8m81
Xpmos_5p04310591302048_3v256x8m81_0 vdd pmos_5p04310591302047_3v256x8m81_0/S vdd pmos_5p04310591302048_3v256x8m81_0/S
+ pmos_5p04310591302048_3v256x8m81
Xpmos_5p04310591302013_3v256x8m81_0 pmos_5p04310591302013_3v256x8m81_0/D se pmos_5p04310591302051_3v256x8m81_0/D
+ se se vdd pmos_5p04310591302013_3v256x8m81
Xnmos_5p04310591302046_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D vss pmos_5p04310591302051_3v256x8m81_0/D
+ pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ q pmos_5p04310591302051_3v256x8m81_0/D vss nmos_5p04310591302046_3v256x8m81
Xpmos_5p04310591302049_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D vdd pmos_5p04310591302051_3v256x8m81_0/D
+ pmos_5p04310591302051_3v256x8m81_0/D q pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ pmos_5p04310591302051_3v256x8m81_0/D vdd pmos_5p04310591302049_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D qp qp vdd
+ pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_1 vdd pmos_5p04310591302048_3v256x8m81_0/S pmos_5p04310591302048_3v256x8m81_0/S
+ vdd pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81
Xpmos_1p2$$171625516_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D vdd vdd pmos_5p04310591302038_3v256x8m81_0/D
+ pmos_5p04310591302013_3v256x8m81_0/D pmos_1p2$$171625516_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D se vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302038_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ vdd vdd pmos_5p04310591302038_3v256x8m81
X0 vss pmos_5p04310591302038_3v256x8m81_0/D pmos_5p04310591302013_3v256x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss se pmos_5p04310591302014_3v256x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X2 pmos_5p04310591302047_3v256x8m81_0/S GWE vss vss nfet_03v3 ad=0.3278p pd=2.37u as=0.3278p ps=2.37u w=0.745u l=0.28u
.ends

.subckt pmos_5p0431059130209_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_5p0431059130207_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt nmos_1p2$$46884908_3v256x8m81 nmos_5p0431059130207_3v256x8m81_0/S a_n14_n34#
+ nmos_5p0431059130207_3v256x8m81_0/D VSUBS
Xnmos_5p0431059130207_3v256x8m81_0 nmos_5p0431059130207_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130207_3v256x8m81_0/S VSUBS nmos_5p0431059130207_3v256x8m81
.ends

.subckt pmos_5p0431059130201_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt pmos_1p2$$46889004_3v256x8m81 pmos_5p0431059130201_3v256x8m81_0/D a_n14_n34#
+ pmos_5p0431059130201_3v256x8m81_0/S w_n133_n66#
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v256x8m81_0/S pmos_5p0431059130201_3v256x8m81
.ends

.subckt nmos_5p0431059130205_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_1p2$$46883884_3v256x8m81 nmos_5p0431059130205_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130205_3v256x8m81_0 nmos_5p0431059130205_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v256x8m81_0/S VSUBS nmos_5p0431059130205_3v256x8m81
.ends

.subckt pmos_5p0431059130206_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302010_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46273580_3v256x8m81 w_n133_n66# a_n42_n34# pmos_5p0431059130203_3v256x8m81_0/S
+ a_118_n34# pmos_5p0431059130203_3v256x8m81_0/D
Xpmos_5p0431059130203_3v256x8m81_0 pmos_5p0431059130203_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p0431059130203_3v256x8m81_0/S pmos_5p0431059130203_3v256x8m81
.ends

.subckt nmos_5p04310591302011_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt pmos_1p2$$46885932_3v256x8m81 pmos_5p0431059130206_3v256x8m81_0/S pmos_5p0431059130206_3v256x8m81_0/D
+ a_118_89# a_n42_89# w_n133_n65#
Xpmos_5p0431059130206_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D a_n42_89# a_118_89#
+ w_n133_n65# pmos_5p0431059130206_3v256x8m81_0/S pmos_5p0431059130206_3v256x8m81
.ends

.subckt nmos_1p2$$46563372_3v256x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt pmos_5p0431059130204_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt pmos_1p2$$46887980_3v256x8m81 w_n133_n66# pmos_5p0431059130204_3v256x8m81_0/S
+ a_n14_n34# pmos_5p0431059130204_3v256x8m81_0/D
Xpmos_5p0431059130204_3v256x8m81_0 pmos_5p0431059130204_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130204_3v256x8m81_0/S pmos_5p0431059130204_3v256x8m81
.ends

.subckt din_3v256x8m81 d db datain wep men pmos_5p0431059130206_3v256x8m81_0/D vss
+ vdd m1_114_5647#
Xpmos_5p0431059130209_3v256x8m81_0 vdd pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ vdd pmos_5p0431059130209_3v256x8m81_0/S pmos_5p0431059130209_3v256x8m81
Xnmos_1p2$$46884908_3v256x8m81_0 vss pmos_5p0431059130201_3v256x8m81_0/S pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ vss nmos_1p2$$46884908_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_0 pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ a_357_4344# d vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D nmos_5p04310591302011_3v256x8m81_1/D
+ pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S pmos_5p0431059130201_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_0 pmos_5p0431059130209_3v256x8m81_0/S wep db vss nmos_1p2$$46883884_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_5p0431059130209_3v256x8m81_0/S a_357_4344# db
+ vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130206_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D datain pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130206_3v256x8m81_0/S pmos_5p0431059130206_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_1 vss pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pmos_5p0431059130209_3v256x8m81_0/S vss nmos_1p2$$46883884_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 vss nmos_5p04310591302011_3v256x8m81_1/D pmos_5p0431059130201_3v256x8m81_0/S
+ vss nmos_5p04310591302010_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D men pmos_5p0431059130206_3v256x8m81_0/D
+ men pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D pmos_1p2$$46273580_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_2 pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ wep d vss nmos_1p2$$46883884_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_1 pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_1p2$$46273580_3v256x8m81
Xnmos_5p04310591302011_3v256x8m81_0 vss datain pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81_0/S vss nmos_5p04310591302011_3v256x8m81
Xnmos_5p04310591302011_3v256x8m81_1 nmos_5p04310591302011_3v256x8m81_1/D pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ men pmos_5p0431059130206_3v256x8m81_0/S vss nmos_5p04310591302011_3v256x8m81
Xpmos_1p2$$46885932_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/S nmos_5p04310591302011_3v256x8m81_1/D
+ pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D men pmos_5p0431059130206_3v256x8m81_0/D
+ pmos_1p2$$46885932_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/S vss pmos_5p0431059130206_3v256x8m81_0/S
+ vss nmos_1p2$$46563372_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_1 men vss pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ vss nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_0 vdd vdd pmos_5p0431059130201_3v256x8m81_0/S pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81
X0 vdd wep a_357_4344# vdd pfet_03v3 ad=0.38572p pd=2.5u as=0.1859p ps=1.23u w=0.695u l=0.28u
X1 a_357_4344# wep vdd vdd pfet_03v3 ad=0.1859p pd=1.23u as=0.38572p ps=2.5u w=0.695u l=0.28u
X2 a_357_4344# wep vss vss nfet_03v3 ad=0.28355p pd=2.13u as=0.3103p ps=2.23u w=0.535u l=0.28u
.ends

.subckt nmos_1p2$$202596396_3v256x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt pmos_5p04310591302041_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt pmos_1p2$$202585132_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n119_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n119_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_5p04310591302043_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
.ends

.subckt nmos_1p2$$202598444_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt pmos_1p2$$202584108_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_1p2$$202587180_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt nmos_5p04310591302039_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302020_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$202586156_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt nmos_1p2$$202595372_3v256x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302042_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# VSUBS
X0 D a_265_n44# S VSUBS nfet_03v3 ad=0.1628p pd=1.62u as=97.125f ps=0.895u w=0.37u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=96.2f pd=0.89u as=0.1628p ps=1.62u w=0.37u l=0.28u
X2 S a_104_n44# D VSUBS nfet_03v3 ad=97.125f pd=0.895u as=96.2f ps=0.89u w=0.37u l=0.28u
.ends

.subckt nmos_1p2$$202594348_3v256x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
.ends

.subckt pmos_1p2$$202583084_3v256x8m81 a_n42_n34# pmos_5p04310591302035_3v256x8m81_0/S
+ w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/D a_118_n34#
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S pmos_5p04310591302035_3v256x8m81
.ends

.subckt wen_wm1_3v256x8m81 GWEN men wep wen vdd vss
Xnmos_1p2$$202596396_3v256x8m81_0 pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ vss pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D vss nmos_1p2$$202596396_3v256x8m81
Xnmos_1p2$$202596396_3v256x8m81_1 pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/D vss vss nmos_1p2$$202596396_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_5/D
+ vdd pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81_0/S vdd vdd pmos_5p04310591302035_3v256x8m81
Xpmos_1p2$$202585132_3v256x8m81_0 vdd pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D vdd pmos_1p2$$202585132_3v256x8m81
Xpmos_5p04310591302043_3v256x8m81_0 wep pmos_5p04310591302035_3v256x8m81_0/D vdd pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_5p04310591302035_3v256x8m81_0/D vdd pmos_5p04310591302043_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 vss pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_5p04310591302020_3v256x8m81_0/S vss nmos_5p04310591302010_3v256x8m81
Xnmos_1p2$$202598444_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81_5/D
+ pmos_5p04310591302014_3v256x8m81_1/D vss nmos_1p2$$202598444_3v256x8m81
Xpmos_1p2$$202584108_3v256x8m81_0 pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S vdd vdd pmos_1p2$$202584108_3v256x8m81
Xpmos_1p2$$202587180_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_4/D
+ pmos_5p04310591302041_3v256x8m81_0/S vdd pmos_1p2$$202587180_3v256x8m81
Xnmos_5p04310591302039_3v256x8m81_0 men pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S
+ vss nmos_5p04310591302039_3v256x8m81
Xpmos_5p04310591302020_3v256x8m81_0 men pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D vdd pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81
Xpmos_1p2$$202586156_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ vdd vdd pmos_1p2$$202586156_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/D vss nmos_1p2$$202595372_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_1 pmos_5p04310591302041_3v256x8m81_0/S pmos_1p2$$202584108_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/S
+ vss vss nmos_1p2$$202595372_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_2/S wen vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xnmos_5p04310591302042_3v256x8m81_0 wep pmos_5p04310591302035_3v256x8m81_0/D vss pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_5p04310591302035_3v256x8m81_0/D vss nmos_5p04310591302042_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_1 pmos_5p04310591302014_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_2/D
+ vdd vdd pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_2 pmos_5p04310591302014_3v256x8m81_2/D GWEN vdd
+ pmos_5p04310591302014_3v256x8m81_2/S pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_3 pmos_5p04310591302014_3v256x8m81_5/S men vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xnmos_1p2$$202594348_3v256x8m81_0 pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D vss vss nmos_1p2$$202594348_3v256x8m81
Xpmos_1p2$$202583084_3v256x8m81_0 pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ vdd vdd pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_1p2$$202585132_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_1p2$$202583084_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_4 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302014_3v256x8m81_5/D
+ vdd vdd pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_5 pmos_5p04310591302014_3v256x8m81_5/D vss vdd pmos_5p04310591302014_3v256x8m81_5/S
+ pmos_5p04310591302014_3v256x8m81
X0 pmos_5p04310591302014_3v256x8m81_5/D men vss vss nfet_03v3 ad=0.1651p pd=1.155u as=0.2794p ps=2.15u w=0.635u l=0.28u
X1 vss GWEN pmos_5p04310591302014_3v256x8m81_2/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
X2 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302014_3v256x8m81_5/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X3 pmos_5p04310591302014_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_2/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X4 vss vss pmos_5p04310591302014_3v256x8m81_5/D vss nfet_03v3 ad=0.2794p pd=2.15u as=0.1651p ps=1.155u w=0.635u l=0.28u
X5 pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S vss vss nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
X6 pmos_5p04310591302014_3v256x8m81_2/D wen vss vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p0431059130200_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt nmos_1p2$$47119404_3v256x8m81 nmos_5p0431059130200_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130200_3v256x8m81_0 nmos_5p0431059130200_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v256x8m81_0/S VSUBS nmos_5p0431059130200_3v256x8m81
.ends

.subckt nmos_5p0431059130202_3v256x8m81 D a_n32_n44# a_136_n44# S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=91.3f pd=0.92u as=0.1561p ps=1.64u w=0.265u l=0.28u
X1 S a_136_n44# D VSUBS nfet_03v3 ad=0.15742p pd=1.65u as=91.3f ps=0.92u w=0.265u l=0.28u
.ends

.subckt ypass_gate_3v256x8m81 vss b bb ypass pcb m3_n41_6881# m3_n41_5924# m3_n41_6639#
+ m3_n41_4610# pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ m3_n41_5682# a_94_7110# vdd m3_n41_5198# m3_n41_5440# m3_n41_6156# via1_2_3v256x8m81_0/VSUBS
+ db
Xnmos_1p2$$47119404_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass b via1_2_3v256x8m81_0/VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_1p2$$47119404_3v256x8m81_3 db ypass bb via1_2_3v256x8m81_0/VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D ypass ypass
+ via1_2_3v256x8m81_0/VSUBS via1_2_3v256x8m81_0/VSUBS nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 b pcb vdd bb pmos_5p0431059130201_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ nmos_5p0431059130202_3v256x8m81_0/D b vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 db nmos_5p0431059130202_3v256x8m81_0/D vdd bb pmos_5p0431059130201_3v256x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.92722p pd=4.34u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 b pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.93515p ps=4.35u w=1.585u l=0.28u
X2 nmos_5p0431059130202_3v256x8m81_0/D ypass vdd vdd pfet_03v3 ad=0.26235p pd=1.45u as=0.46218p ps=2.72u w=0.695u l=0.28u
X3 vdd ypass nmos_5p0431059130202_3v256x8m81_0/D vdd pfet_03v3 ad=0.39963p pd=2.54u as=0.26235p ps=1.45u w=0.695u l=0.28u
X4 vdd pcb bb vdd pfet_03v3 ad=0.93015p pd=4.35u as=0.4134p ps=2.11u w=1.59u l=0.28u
X5 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=0.9381p ps=4.36u w=1.59u l=0.28u
.ends

.subckt ypass_gate_a_3v256x8m81 vss b bb ypass pcb m3_n41_6881# a_64_7110# m3_n41_5924#
+ m3_n41_6639# m3_n41_4610# pmos_5p0431059130201_3v256x8m81_0/D m3_n41_5682# via1_2_3v256x8m81_0/VSUBS
+ vdd pmos_5p0431059130201_3v256x8m81_1/D pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ m3_n41_5198# m3_n41_5440# m3_n41_6156#
Xnmos_1p2$$47119404_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass pmos_5p0431059130201_3v256x8m81_0/D via1_2_3v256x8m81_0/VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_1p2$$47119404_3v256x8m81_3 pmos_5p0431059130201_3v256x8m81_1/D ypass bb via1_2_3v256x8m81_0/VSUBS
+ nmos_1p2$$47119404_3v256x8m81
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D ypass ypass
+ via1_2_3v256x8m81_0/VSUBS via1_2_3v256x8m81_0/VSUBS nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D pcb vdd bb
+ pmos_5p0431059130201_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ nmos_5p0431059130202_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/D vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 pmos_5p0431059130201_3v256x8m81_1/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v256x8m81
X0 vdd pcb pmos_5p0431059130201_3v256x8m81_0/D vdd pfet_03v3 ad=1.06988p pd=4.52u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 pmos_5p0431059130201_3v256x8m81_0/D pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.99855p ps=4.43u w=1.585u l=0.28u
X2 vdd ypass nmos_5p0431059130202_3v256x8m81_0/D vdd pfet_03v3 ad=0.5143p pd=2.87u as=0.34055p ps=1.675u w=0.695u l=0.28u
X3 vdd pcb bb vdd pfet_03v3 ad=1.07325p pd=4.53u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=1.0017p ps=4.44u w=1.59u l=0.28u
X5 nmos_5p0431059130202_3v256x8m81_0/D ypass vdd vdd pfet_03v3 ad=0.34055p pd=1.675u as=0.38572p ps=2.5u w=0.695u l=0.28u
.ends

.subckt mux821_3v256x8m81 ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_6/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_6/b ypass_gate_a_3v256x8m81_0/ypass ypass_gate_3v256x8m81_7/bb
+ ypass_gate_3v256x8m81_4/bb ypass_gate_3v256x8m81_1/bb ypass_gate_3v256x8m81_1/b
+ ypass_gate_3v256x8m81_1/db ypass_gate_3v256x8m81_1/ypass ypass_gate_3v256x8m81_4/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_3/b ypass_gate_3v256x8m81_2/ypass ypass_gate_3v256x8m81_3/ypass
+ ypass_gate_3v256x8m81_4/ypass ypass_gate_3v256x8m81_5/b ypass_gate_3v256x8m81_5/ypass
+ ypass_gate_3v256x8m81_6/ypass ypass_gate_3v256x8m81_7/ypass ypass_gate_3v256x8m81_7/b
+ ypass_gate_3v256x8m81_6/bb ypass_gate_3v256x8m81_3/bb ypass_gate_3v256x8m81_7/db
+ ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81_5/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_a_3v256x8m81_0/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_a_3v256x8m81_0/bb ypass_gate_3v256x8m81_2/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_2/b
+ ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_7/m3_n41_6156#
+ ypass_gate_3v256x8m81_5/bb ypass_gate_3v256x8m81_2/bb ypass_gate_3v256x8m81_4/b
+ ypass_gate_3v256x8m81_3/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_1/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_4/db VSUBS ypass_gate_3v256x8m81_7/m3_n41_6881#
Xypass_gate_3v256x8m81_1 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_1/b ypass_gate_3v256x8m81_1/bb
+ ypass_gate_3v256x8m81_1/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_1/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_1/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_2 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_2/b ypass_gate_3v256x8m81_2/bb
+ ypass_gate_3v256x8m81_2/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_2/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_4/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_3 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_3/b ypass_gate_3v256x8m81_3/bb
+ ypass_gate_3v256x8m81_3/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_3/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_4 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_4/b ypass_gate_3v256x8m81_4/bb
+ ypass_gate_3v256x8m81_4/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_4/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_4/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_5 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_5/b ypass_gate_3v256x8m81_5/bb
+ ypass_gate_3v256x8m81_5/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_5/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_6 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_6/b ypass_gate_3v256x8m81_6/bb
+ ypass_gate_3v256x8m81_6/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_6/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_7/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_7 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/b ypass_gate_3v256x8m81_7/bb
+ ypass_gate_3v256x8m81_7/ypass ypass_gate_3v256x8m81_7/pcb ypass_gate_3v256x8m81_7/m3_n41_6881#
+ ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/vdd
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v256x8m81_7/db ypass_gate_3v256x8m81
Xypass_gate_a_3v256x8m81_0 ypass_gate_3v256x8m81_7/vss ypass_gate_a_3v256x8m81_0/b
+ ypass_gate_a_3v256x8m81_0/bb ypass_gate_a_3v256x8m81_0/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/a_94_7110# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# VSUBS ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_1/db
+ ypass_gate_a_3v256x8m81_0/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ ypass_gate_a_3v256x8m81
.ends

.subckt pmos_5p04310591302018_3v256x8m81 a_20_n45# D a_181_n45# a_502_n45# a_662_n45#
+ a_n140_n45# S a_341_n45# w_n314_n86#
X0 S a_341_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_662_n45# D w_n314_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_502_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 S a_20_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_181_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X5 D a_n140_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46549036_3v256x8m81 a_327_n34# w_n188_n50# pmos_5p04310591302018_3v256x8m81_0/S
+ a_488_n34# a_n154_n34# a_167_n34# pmos_5p04310591302018_3v256x8m81_0/D a_6_n34#
+ a_648_n34#
Xpmos_5p04310591302018_3v256x8m81_0 a_6_n34# pmos_5p04310591302018_3v256x8m81_0/D
+ a_167_n34# a_488_n34# a_648_n34# a_n154_n34# pmos_5p04310591302018_3v256x8m81_0/S
+ a_327_n34# w_n188_n50# pmos_5p04310591302018_3v256x8m81
.ends

.subckt pmos_5p04310591302021_3v256x8m81 a_76_n44# D a_n84_n44# w_n258_n86# S a_237_n44#
+ a_397_n44#
X0 S a_397_n44# D w_n258_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1092p ps=0.94u w=0.42u l=0.28u
X1 D a_237_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.11025p ps=0.945u w=0.42u l=0.28u
X2 D a_n84_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.1848p ps=1.72u w=0.42u l=0.28u
X3 S a_76_n44# D w_n258_n86# pfet_03v3 ad=0.11025p pd=0.945u as=0.1092p ps=0.94u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46896172_3v256x8m81 w_n133_n66# pmos_5p04310591302021_3v256x8m81_0/S
+ pmos_5p04310591302021_3v256x8m81_0/a_n84_n44# pmos_5p04310591302021_3v256x8m81_0/D
+ pmos_5p04310591302021_3v256x8m81_0/a_76_n44# pmos_5p04310591302021_3v256x8m81_0/a_237_n44#
+ pmos_5p04310591302021_3v256x8m81_0/a_397_n44#
Xpmos_5p04310591302021_3v256x8m81_0 pmos_5p04310591302021_3v256x8m81_0/a_76_n44# pmos_5p04310591302021_3v256x8m81_0/D
+ pmos_5p04310591302021_3v256x8m81_0/a_n84_n44# w_n133_n66# pmos_5p04310591302021_3v256x8m81_0/S
+ pmos_5p04310591302021_3v256x8m81_0/a_237_n44# pmos_5p04310591302021_3v256x8m81_0/a_397_n44#
+ pmos_5p04310591302021_3v256x8m81
.ends

.subckt pmos_1p2$$46897196_3v256x8m81 w_n133_n66# a_n42_n34# pmos_5p04310591302020_3v256x8m81_0/D
+ a_118_n34# pmos_5p04310591302020_3v256x8m81_0/S
Xpmos_5p04310591302020_3v256x8m81_0 pmos_5p04310591302020_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302020_3v256x8m81_0/S pmos_5p04310591302020_3v256x8m81
.ends

.subckt nmos_5p04310591302015_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6996p pd=4.06u as=0.6996p ps=4.06u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46553132_3v256x8m81 nmos_5p04310591302015_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302015_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302015_3v256x8m81_0 nmos_5p04310591302015_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302015_3v256x8m81_0/S VSUBS nmos_5p04310591302015_3v256x8m81
.ends

.subckt nmos_1p2$$45107244_3v256x8m81 a_223_n34# a_383_n34# nmos_5p04310591302012_3v256x8m81_0/S
+ a_n96_n34# a_63_n34# nmos_5p04310591302012_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302012_3v256x8m81_0 a_n96_n34# nmos_5p04310591302012_3v256x8m81_0/D
+ a_63_n34# nmos_5p04310591302012_3v256x8m81_0/S a_223_n34# a_383_n34# VSUBS nmos_5p04310591302012_3v256x8m81
.ends

.subckt nmos_5p04310591302016_3v256x8m81 a_124_n45# a_284_n45# D a_446_n45# a_768_n45#
+ a_n198_n45# a_n38_n45# a_606_n45# S a_928_n45# VSUBS
X0 S a_928_n45# D VSUBS nfet_03v3 ad=0.7155p pd=4.08u as=0.4134p ps=2.11u w=1.59u l=0.28u
X1 D a_n198_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.70755p ps=4.07u w=1.59u l=0.28u
X2 S a_n38_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X3 S a_606_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 D a_768_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X5 D a_446_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X6 S a_284_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X7 D a_124_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46552108_3v256x8m81 nmos_5p04310591302016_3v256x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_284_n45# nmos_5p04310591302016_3v256x8m81_0/a_446_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_768_n45# nmos_5p04310591302016_3v256x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v256x8m81_0/S nmos_5p04310591302016_3v256x8m81_0/a_n198_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_606_n45# nmos_5p04310591302016_3v256x8m81_0/a_928_n45#
+ nmos_5p04310591302016_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302016_3v256x8m81_0 nmos_5p04310591302016_3v256x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_284_n45# nmos_5p04310591302016_3v256x8m81_0/D
+ nmos_5p04310591302016_3v256x8m81_0/a_446_n45# nmos_5p04310591302016_3v256x8m81_0/a_768_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_n198_n45# nmos_5p04310591302016_3v256x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_606_n45# nmos_5p04310591302016_3v256x8m81_0/S
+ nmos_5p04310591302016_3v256x8m81_0/a_928_n45# VSUBS nmos_5p04310591302016_3v256x8m81
.ends

.subckt pmos_5p04310591302019_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46898220_3v256x8m81 w_n133_n66# a_n14_84# pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_5p04310591302019_3v256x8m81_0/D
Xpmos_5p04310591302019_3v256x8m81_0 pmos_5p04310591302019_3v256x8m81_0/D a_n14_84#
+ w_n133_n66# pmos_5p04310591302019_3v256x8m81_0/S pmos_5p04310591302019_3v256x8m81
.ends

.subckt nmos_5p04310591302017_3v256x8m81 a_n37_n44# D a_929_n44# a_125_n44# a_285_n44#
+ a_447_n44# a_769_n44# S a_607_n44# a_n197_n44# VSUBS
X0 D a_769_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X1 D a_447_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X2 D a_n197_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X3 S a_n37_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X4 S a_285_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X5 D a_125_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X6 S a_929_n44# D VSUBS nfet_03v3 ad=0.58963p pd=3.54u as=0.3445p ps=1.845u w=1.325u l=0.28u
X7 S a_607_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_1p2$$46550060_3v256x8m81 nmos_5p04310591302017_3v256x8m81_0/D a_915_n34#
+ a_111_n34# a_271_n34# a_433_n34# a_593_n34# a_n51_n34# a_755_n34# a_n210_n34# nmos_5p04310591302017_3v256x8m81_0/S
+ VSUBS
Xnmos_5p04310591302017_3v256x8m81_0 a_n51_n34# nmos_5p04310591302017_3v256x8m81_0/D
+ a_915_n34# a_111_n34# a_271_n34# a_433_n34# a_755_n34# nmos_5p04310591302017_3v256x8m81_0/S
+ a_593_n34# a_n210_n34# VSUBS nmos_5p04310591302017_3v256x8m81
.ends

.subckt nmos_1p2$$46551084_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt sa_3v256x8m81 qp wep se pcb d vdd vss
Xpmos_1p2$$46549036_3v256x8m81_0 qp vdd vdd pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S qp qp pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46549036_3v256x8m81
Xpmos_1p2$$46896172_3v256x8m81_0 d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46896172_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_0 d se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ se d pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_1 d se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ se d pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_2 d se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ se d pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_3 d se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ se d pmos_1p2$$46897196_3v256x8m81
Xnmos_1p2$$46553132_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_3v256x8m81
Xnmos_1p2$$46553132_3v256x8m81_1 vss vss pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ vss nmos_1p2$$46553132_3v256x8m81
Xnmos_1p2$$45107244_3v256x8m81_0 qp qp qp pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ qp vss vss nmos_1p2$$45107244_3v256x8m81
Xnmos_1p2$$46552108_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D vss nmos_1p2$$46552108_3v256x8m81
Xpmos_1p2$$46898220_3v256x8m81_0 d d d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81
Xnmos_1p2$$46550060_3v256x8m81_0 nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ se se se se se se se se vss vss nmos_1p2$$46550060_3v256x8m81
Xpmos_1p2$$46898220_3v256x8m81_1 d d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ d pmos_1p2$$46898220_3v256x8m81
Xpmos_1p2$$46286892_3v256x8m81_0 d d pcb pcb pcb d pmos_1p2$$46286892_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 vss pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ qp vss nmos_1p2$$46551084_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pcb pmos_1p2$$46285868_3v256x8m81
.ends

.subckt saout_R_m2_3v256x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWE GWEN
+ datain b[5] b[4] b[2] b[1] b[0] bb[6] q bb[3] bb[0] bb[1] pcb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ bb[5] sa_3v256x8m81_0/pcb WEN mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b bb[2]
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb b[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass
+ din_3v256x8m81_0/men mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass bb[4] b[6]
+ ypass[7] m2_26_12231# mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ bb[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ vss vdd
Xsacntl_2_3v256x8m81_0 sa_3v256x8m81_0/pcb sa_3v256x8m81_0/se din_3v256x8m81_0/men
+ sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_1/S sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_2/S
+ vss vdd sacntl_2_3v256x8m81
Xoutbuf_oe_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qp sa_3v256x8m81_0/se q
+ GWE vss vdd outbuf_oe_3v256x8m81
Xdin_3v256x8m81_0 vdd vdd datain sa_3v256x8m81_0/wep din_3v256x8m81_0/men vdd vss
+ vdd sa_3v256x8m81_0/pcb din_3v256x8m81
Xwen_wm1_3v256x8m81_0 GWEN din_3v256x8m81_0/men sa_3v256x8m81_0/wep WEN vdd vss wen_wm1_3v256x8m81
Xmux821_3v256x8m81_0 mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb bb[5] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ b[6] vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass vdd vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass
+ ypass[7] b[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb bb[2] vdd vdd vdd vdd bb[7] vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass sa_3v256x8m81_0/pcb ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b m2_26_12231# vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb bb[4] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass
+ vdd vss mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81
Xsa_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/wep sa_3v256x8m81_0/se sa_3v256x8m81_0/pcb
+ vdd vdd vss sa_3v256x8m81
.ends

.subckt x018SRAM_cell1_2x_3v256x8m81 018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_3v256x8m81_0/a_62_178# 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_62_178# VSUBS
X018SRAM_cell1_3v256x8m81_0 018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_3v256x8m81_0/a_62_178# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_62_178# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v256x8m81
.ends

.subckt Cell_array8x8_3v256x8m81 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS
X018SRAM_cell1_2x_3v256x8m81_0[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
.ends

.subckt saout_m2_3v256x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWEN GWE
+ bb[1] bb[4] bb[7] bb[6] b[5] b[7] b[2] q pcb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ b[6] bb[2] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass WEN mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb bb[5] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ b[4] din_3v256x8m81_0/men mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b outbuf_oe_3v256x8m81_0/GWE
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[3] b[1] ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass b[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass vss mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass vdd
Xsacntl_2_3v256x8m81_0 pcb sa_3v256x8m81_0/se din_3v256x8m81_0/men sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_1/S
+ sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_2/S vss vdd sacntl_2_3v256x8m81
Xoutbuf_oe_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qp sa_3v256x8m81_0/se q
+ outbuf_oe_3v256x8m81_0/GWE vss vdd outbuf_oe_3v256x8m81
Xdin_3v256x8m81_0 vdd vdd vdd sa_3v256x8m81_0/wep din_3v256x8m81_0/men vdd vss vdd
+ pcb din_3v256x8m81
Xwen_wm1_3v256x8m81_0 GWEN din_3v256x8m81_0/men sa_3v256x8m81_0/wep WEN vdd vss wen_wm1_3v256x8m81
Xmux821_3v256x8m81_0 mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ vdd b[6] mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ bb[2] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb b[1] vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ vdd vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass b[4] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[5] vdd vdd vdd vdd mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb vdd mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass pcb ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ b[3] vss vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ bb[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass vdd vss mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81
Xsa_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/wep sa_3v256x8m81_0/se pcb vdd
+ vdd vss sa_3v256x8m81
.ends

.subckt col_256a_3v256x8m81 ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] ypass[7]
+ GWE WL[32] WL[31] WL[30] WL[20] WL[11] WL[10] WL[7] WL[18] WL[17] WL[16] WL[15]
+ WL[14] WL[13] WL[27] WL[26] ypass[6] ypass[2] b[1] b[7] b[10] b[13] b[16] b[22]
+ b[28] din[1] din[3] din[2] din[0] q[0] q[1] q[2] q[3] b[29] b[23] b[20] b[14] b[11]
+ b[8] bb[0] bb[1] bb[2] bb[8] bb[9] bb[11] bb[12] bb[13] bb[14] bb[15] bb[19] bb[21]
+ bb[22] bb[24] bb[26] bb[28] bb[29] bb[30] bb[31] b[30] b[27] b[0] b[3] b[18] pcb[0]
+ pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1] WEN[0] saout_R_m2_3v256x8m81_0/q saout_R_m2_3v256x8m81_1/datain
+ saout_m2_3v256x8m81_4/GWEN WL[1] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_4/q WL[4] men saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[21] m3_n771_22409# saout_R_m2_3v256x8m81_0/datain b[9] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[24] saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_0/GWE saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b b[25] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb WL[5] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_4/GWE saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[8] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/b[1]
+ saout_R_m2_3v256x8m81_1/bb[5] WL[25] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_4/b[6] saout_m2_3v256x8m81_3/bb[5] WL[2] WL[28] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_0/b[3] saout_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_1/q
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/q WL[22] saout_m2_3v256x8m81_4/b[3] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ b[31] saout_R_m2_3v256x8m81_1/GWE saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[9] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb bb[4]
+ WL[12] b[12] saout_m2_3v256x8m81_4/bb[5] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[3] saout_m2_3v256x8m81_3/b[4] WL[29] b[5] WL[6] saout_R_m2_3v256x8m81_0/bb[4]
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_1/b[3]
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb bb[17] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/b[6] saout_R_m2_3v256x8m81_1/bb[4] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_0/bb[2] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/b[3] WL[23] saout_R_m2_3v256x8m81_1/bb[7] bb[10] WL[19] VSS
+ VDD WL[0] bb[6]
Xsaout_R_m2_3v256x8m81_0 saout_R_m2_3v256x8m81_0/ypass[2] saout_R_m2_3v256x8m81_0/ypass[3]
+ saout_R_m2_3v256x8m81_0/ypass[4] saout_R_m2_3v256x8m81_0/ypass[5] saout_R_m2_3v256x8m81_0/ypass[6]
+ saout_R_m2_3v256x8m81_0/GWE saout_m2_3v256x8m81_4/GWEN saout_R_m2_3v256x8m81_0/datain
+ saout_R_m2_3v256x8m81_0/b[5] saout_R_m2_3v256x8m81_0/b[4] saout_R_m2_3v256x8m81_0/b[2]
+ saout_R_m2_3v256x8m81_0/b[1] saout_R_m2_3v256x8m81_0/b[0] saout_R_m2_3v256x8m81_0/bb[6]
+ saout_R_m2_3v256x8m81_0/q saout_R_m2_3v256x8m81_0/bb[3] saout_R_m2_3v256x8m81_0/bb[0]
+ saout_R_m2_3v256x8m81_0/bb[1] saout_R_m2_3v256x8m81_0/pcb saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ bb[4] saout_R_m2_3v256x8m81_0/sa_3v256x8m81_0/pcb WEN[0] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_0/bb[2] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_0/b[3] ypass[2] men ypass[0] saout_R_m2_3v256x8m81_0/bb[4]
+ b[5] ypass[5] VSS ypass[1] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b ypass[4] bb[6]
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb ypass[6]
+ ypass[3] ypass[7] VSS VDD saout_R_m2_3v256x8m81
Xsaout_R_m2_3v256x8m81_1 saout_R_m2_3v256x8m81_1/ypass[2] saout_R_m2_3v256x8m81_1/ypass[3]
+ saout_R_m2_3v256x8m81_1/ypass[4] saout_R_m2_3v256x8m81_1/ypass[5] saout_R_m2_3v256x8m81_1/ypass[6]
+ saout_R_m2_3v256x8m81_1/GWE saout_m2_3v256x8m81_4/GWEN saout_R_m2_3v256x8m81_1/datain
+ saout_R_m2_3v256x8m81_1/b[5] saout_R_m2_3v256x8m81_1/b[4] saout_R_m2_3v256x8m81_1/b[2]
+ saout_R_m2_3v256x8m81_1/b[1] saout_R_m2_3v256x8m81_1/b[0] saout_R_m2_3v256x8m81_1/bb[6]
+ saout_R_m2_3v256x8m81_1/q saout_R_m2_3v256x8m81_1/bb[3] saout_R_m2_3v256x8m81_1/bb[0]
+ saout_R_m2_3v256x8m81_1/bb[1] saout_R_m2_3v256x8m81_1/pcb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb WEN[2]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b b[18] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_1/b[3] ypass[2] men ypass[0] saout_R_m2_3v256x8m81_1/bb[4]
+ saout_R_m2_3v256x8m81_1/b[6] ypass[5] VSS ypass[1] bb[17] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ ypass[4] saout_R_m2_3v256x8m81_1/bb[7] b[16] ypass[6] ypass[3] ypass[7] VSS VDD
+ saout_R_m2_3v256x8m81
XCell_array8x8_3v256x8m81_0 saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b bb[8] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ b[10] saout_R_m2_3v256x8m81_0/b[3] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[6] b[9] b[29] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb WL[22] bb[11]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_0/bb[4]
+ b[25] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_1/bb[4]
+ bb[10] bb[30] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_3/b[1] WL[28] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[23] b[12] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[29] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b b[18] saout_m2_3v256x8m81_4/b[3]
+ b[31] b[16] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_1/b[6]
+ WL[24] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_m2_3v256x8m81_4/bb[5]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[4] WL[10] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ WL[8] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb WL[17]
+ saout_R_m2_3v256x8m81_1/b[3] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[0] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[19] bb[17] bb[4] WL[9] WL[3] WL[6] saout_R_m2_3v256x8m81_0/bb[2] saout_m2_3v256x8m81_3/b[3]
+ WL[16] saout_m2_3v256x8m81_3/b[6] WL[1] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[11] WL[21] saout_R_m2_3v256x8m81_1/bb[7] WL[31] WL[2] bb[24] saout_R_m2_3v256x8m81_1/bb[5]
+ WL[20] WL[12] WL[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[5] WL[27] WL[25] WL[26] b[5] WL[30] WL[18] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[15] WL[13] WL[4] saout_m2_3v256x8m81_4/b[6] VDD saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ WL[14] VSS Cell_array8x8_3v256x8m81
Xsaout_m2_3v256x8m81_3 saout_m2_3v256x8m81_3/ypass[2] saout_m2_3v256x8m81_3/ypass[3]
+ saout_m2_3v256x8m81_3/ypass[4] saout_m2_3v256x8m81_3/ypass[5] saout_m2_3v256x8m81_3/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN GWE saout_m2_3v256x8m81_3/bb[1] saout_m2_3v256x8m81_3/bb[4]
+ saout_m2_3v256x8m81_3/bb[7] saout_m2_3v256x8m81_3/bb[6] saout_m2_3v256x8m81_3/b[5]
+ saout_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[2] saout_m2_3v256x8m81_3/q saout_m2_3v256x8m81_3/pcb
+ b[29] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/bb[2] ypass[2] WEN[3] b[31] bb[24]
+ saout_m2_3v256x8m81_3/bb[5] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_3/b[4] men b[25] GWE ypass[0] bb[30] saout_m2_3v256x8m81_3/bb[3]
+ saout_m2_3v256x8m81_3/b[1] ypass[5] ypass[1] saout_m2_3v256x8m81_3/b[3] ypass[4]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ ypass[3] VSS ypass[7] ypass[6] VDD saout_m2_3v256x8m81
Xsaout_m2_3v256x8m81_4 saout_m2_3v256x8m81_4/ypass[2] saout_m2_3v256x8m81_4/ypass[3]
+ saout_m2_3v256x8m81_4/ypass[4] saout_m2_3v256x8m81_4/ypass[5] saout_m2_3v256x8m81_4/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN saout_m2_3v256x8m81_4/GWE saout_m2_3v256x8m81_4/bb[1]
+ saout_m2_3v256x8m81_4/bb[4] saout_m2_3v256x8m81_4/bb[7] saout_m2_3v256x8m81_4/bb[6]
+ saout_m2_3v256x8m81_4/b[5] saout_m2_3v256x8m81_4/b[7] saout_m2_3v256x8m81_4/b[2]
+ saout_m2_3v256x8m81_4/q saout_m2_3v256x8m81_4/pcb saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_4/b[6] bb[10] ypass[2] WEN[1] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb saout_m2_3v256x8m81_4/bb[5]
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb b[12] men b[10]
+ saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE ypass[0] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[11] b[9] ypass[5] ypass[1] saout_m2_3v256x8m81_4/b[3] ypass[4] bb[8] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ ypass[3] VSS ypass[7] ypass[6] VDD saout_m2_3v256x8m81
.ends

.subckt dcap_103_novia_3v256x8m81 w_n205_0# a_n30_42# a_n119_86#
X0 a_n119_86# a_n30_42# a_n119_86# w_n205_0# pfet_03v3 ad=0.4717p pd=3.01u as=0 ps=0 w=1.06u l=1.74u
.ends

.subckt lcol4_256_3v256x8m81 WL[20] WL[19] WL[18] WL[16] WL[14] WL[13] WL[12] WL[10]
+ WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[31] din[1] din[3] din[2]
+ q[1] q[2] q[3] pcb[2] pcb[3] pcb[0] pcb[1] WEN[3] WEN[2] WEN[1] WEN[0] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/GWE
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/q col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/q
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWEN col_256a_3v256x8m81_0/WL[6] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE
+ col_256a_3v256x8m81_0/WL[8] col_256a_3v256x8m81_0/WL[21] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/datain
+ WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/datain
+ WL[27] WL[28] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/q col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/q
+ col_256a_3v256x8m81_0/ypass[0] col_256a_3v256x8m81_0/ypass[1] col_256a_3v256x8m81_0/ypass[2]
+ col_256a_3v256x8m81_0/ypass[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/GWE
+ col_256a_3v256x8m81_0/ypass[4] col_256a_3v256x8m81_0/men col_256a_3v256x8m81_0/WL[10]
+ col_256a_3v256x8m81_0/ypass[5] col_256a_3v256x8m81_0/ypass[6] WL[11] col_256a_3v256x8m81_0/ypass[7]
+ col_256a_3v256x8m81_0/WL[12] col_256a_3v256x8m81_0/GWE WL[29] col_256a_3v256x8m81_0/WL[13]
+ col_256a_3v256x8m81_0/WL[14] WL[30] col_256a_3v256x8m81_0/WL[15] WL[15] col_256a_3v256x8m81_0/WL[17]
+ WL[17] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWE WL[0] col_256a_3v256x8m81_0/WL[19]
+ VSUBS VDD
Xldummy_3v256x4_3v256x8m81_0 WL[5] VDD VSUBS col_256a_3v256x8m81_0/b[16] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/b[16] VDD col_256a_3v256x8m81_0/bb[10] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/WL[21] VDD WL[25] col_256a_3v256x8m81_0/b[10] col_256a_3v256x8m81_0/b[29]
+ VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5] VDD col_256a_3v256x8m81_0/WL[6]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] VSUBS col_256a_3v256x8m81_0/bb[10]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] col_256a_3v256x8m81_0/b[10] WL[7]
+ WL[3] VDD VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[23] VDD WL[22] VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2]
+ WL[4] VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/b[31] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[9] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/bb[24]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/bb[24] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VDD col_256a_3v256x8m81_0/b[5] WL[21] WL[24] VSUBS VSUBS col_256a_3v256x8m81_0/bb[30]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6] WL[0] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7] col_256a_3v256x8m81_0/bb[6]
+ WL[11] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2] col_256a_3v256x8m81_0/b[25]
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/b[25] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4]
+ VDD VDD WL[19] WL[26] col_256a_3v256x8m81_0/b[31] VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3] WL[2] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/bb[11] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6]
+ col_256a_3v256x8m81_0/WL[13] VSUBS VDD VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ VDD VDD col_256a_3v256x8m81_0/bb[4] WL[17] VSUBS WL[28] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/WL[15] VSUBS VDD col_256a_3v256x8m81_0/b[29] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VDD WL[15] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/b[12] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5]
+ col_256a_3v256x8m81_0/WL[17] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2] VDD col_256a_3v256x8m81_0/WL[14]
+ VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSUBS col_256a_3v256x8m81_0/WL[12] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/bb[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ WL[30] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[29] col_256a_3v256x8m81_0/bb[30] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3]
+ VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/WL[10] VSUBS col_256a_3v256x8m81_0/bb[11] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/b[5] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ VDD VDD col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[27] col_256a_3v256x8m81_0/bb[8] VSUBS col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/WL[8] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4] col_256a_3v256x8m81_0/bb[8]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[1] col_256a_3v256x8m81_0/bb[17] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/bb[17] col_256a_3v256x8m81_0/b[9] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VDD col_256a_3v256x8m81_0/WL[19] VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/b[9] VDD col_256a_3v256x8m81_0/b[12] col_256a_3v256x8m81_0/bb[4]
+ ldummy_3v256x4_3v256x8m81
Xcol_256a_3v256x8m81_0 col_256a_3v256x8m81_0/ypass[0] col_256a_3v256x8m81_0/ypass[1]
+ col_256a_3v256x8m81_0/ypass[3] col_256a_3v256x8m81_0/ypass[4] col_256a_3v256x8m81_0/ypass[5]
+ col_256a_3v256x8m81_0/ypass[7] col_256a_3v256x8m81_0/GWE VSUBS WL[30] WL[29] WL[19]
+ WL[11] col_256a_3v256x8m81_0/WL[10] WL[7] WL[17] col_256a_3v256x8m81_0/WL[17] WL[15]
+ col_256a_3v256x8m81_0/WL[15] col_256a_3v256x8m81_0/WL[14] col_256a_3v256x8m81_0/WL[13]
+ WL[26] WL[25] col_256a_3v256x8m81_0/ypass[6] col_256a_3v256x8m81_0/ypass[2] col_256a_3v256x8m81_0/b[1]
+ col_256a_3v256x8m81_0/b[7] col_256a_3v256x8m81_0/b[10] col_256a_3v256x8m81_0/b[13]
+ col_256a_3v256x8m81_0/b[16] col_256a_3v256x8m81_0/b[22] col_256a_3v256x8m81_0/b[28]
+ col_256a_3v256x8m81_0/din[1] col_256a_3v256x8m81_0/din[3] col_256a_3v256x8m81_0/din[2]
+ col_256a_3v256x8m81_0/din[0] col_256a_3v256x8m81_0/q[0] col_256a_3v256x8m81_0/q[1]
+ col_256a_3v256x8m81_0/q[2] col_256a_3v256x8m81_0/q[3] col_256a_3v256x8m81_0/b[29]
+ col_256a_3v256x8m81_0/b[23] col_256a_3v256x8m81_0/b[20] col_256a_3v256x8m81_0/b[14]
+ col_256a_3v256x8m81_0/b[11] col_256a_3v256x8m81_0/b[8] col_256a_3v256x8m81_0/bb[0]
+ col_256a_3v256x8m81_0/bb[1] col_256a_3v256x8m81_0/bb[2] col_256a_3v256x8m81_0/bb[8]
+ col_256a_3v256x8m81_0/bb[9] col_256a_3v256x8m81_0/bb[11] col_256a_3v256x8m81_0/bb[12]
+ col_256a_3v256x8m81_0/bb[13] col_256a_3v256x8m81_0/bb[14] col_256a_3v256x8m81_0/bb[15]
+ col_256a_3v256x8m81_0/bb[19] col_256a_3v256x8m81_0/bb[21] col_256a_3v256x8m81_0/bb[22]
+ col_256a_3v256x8m81_0/bb[24] col_256a_3v256x8m81_0/bb[26] col_256a_3v256x8m81_0/bb[28]
+ col_256a_3v256x8m81_0/bb[29] col_256a_3v256x8m81_0/bb[30] col_256a_3v256x8m81_0/bb[31]
+ col_256a_3v256x8m81_0/b[30] col_256a_3v256x8m81_0/b[27] col_256a_3v256x8m81_0/b[0]
+ col_256a_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/pcb[0]
+ col_256a_3v256x8m81_0/pcb[1] col_256a_3v256x8m81_0/pcb[3] col_256a_3v256x8m81_0/pcb[2]
+ WEN[3] WEN[2] WEN[1] WEN[0] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/q col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/datain
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWEN WL[1] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/q WL[4] col_256a_3v256x8m81_0/men col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/WL[21] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/datain
+ col_256a_3v256x8m81_0/b[9] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[23] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/GWE col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/b[25] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ WL[5] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWE col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/WL[8] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5]
+ WL[24] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5]
+ WL[2] WL[27] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/q col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/q WL[21] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/b[31] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/GWE col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[9] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/bb[4] col_256a_3v256x8m81_0/WL[12] col_256a_3v256x8m81_0/b[12]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[3] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] WL[28] col_256a_3v256x8m81_0/b[5]
+ col_256a_3v256x8m81_0/WL[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/bb[17] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3] WL[22] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7]
+ col_256a_3v256x8m81_0/bb[10] col_256a_3v256x8m81_0/WL[19] VSUBS VDD WL[0] col_256a_3v256x8m81_0/bb[6]
+ col_256a_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[0] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[1] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[2] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[3] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[4] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[5] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[6] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[7] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[8] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[9] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[10] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[11] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[12] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[13] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[14] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[15] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[16] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[17] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[18] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[19] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[20] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[21] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[22] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[23] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[24] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[25] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[26] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[27] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[28] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[29] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[30] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[31] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[32] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[33] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[34] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[35] VDD VSUBS VDD dcap_103_novia_3v256x8m81
.ends

.subckt rarray4_256_3v256x8m81 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11203# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2719# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_11917# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_8779#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_16765#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3931# m3_n1397_3433# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_2221# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_8281# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_19189#
+ m3_n1397_19687# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_18475#
+ m3_n1397_9991# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_12415# m3_n1397_14839# m3_n1397_15553# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_10705#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_4645#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_13627# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_247# m3_n1397_1507# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_5143#
+ m3_n1397_9493# m3_n1397_17263# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_14341#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# m3_n1397_16051# m3_n1397_7069# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_5857#
+ VSUBS
X018SRAM_cell1_2x_3v256x8m81_456 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_467 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_423 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_412 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_434 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_445 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_478 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_401 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_990 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_7 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_220 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_231 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_297 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_286 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_253 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_275 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_242 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_264 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_19 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_457 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_424 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_413 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_468 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_435 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_446 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_479 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_402 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_980 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_8 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_221 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_210 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_298 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_287 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_254 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_276 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_243 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_265 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_232 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1020 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_425 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_414 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_469 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_447 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_458 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_436 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_403 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_9 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_992 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_970 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_200 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_222 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_211 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1010 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_299 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_288 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_255 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_277 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_244 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_266 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_233 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_448 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_426 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_415 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_437 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_459 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_404 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_982 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_960 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_201 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_234 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_223 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1000 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_245 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1022 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_212 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_278 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_289 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_267 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_449 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_416 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_438 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_405 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_427 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_994 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_972 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1012 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_235 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_202 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_257 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_279 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_246 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_268 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_224 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_213 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_439 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_417 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_406 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_428 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_984 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_962 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1002 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_203 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_258 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_269 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_247 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_214 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_225 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_236 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_418 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_429 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_407 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_996 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_974 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_204 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_226 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1014 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_259 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_248 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_215 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_237 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_419 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_408 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_986 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_964 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_216 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_205 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_227 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_238 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1004 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_249 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_409 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_998 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_976 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_217 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_206 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_239 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_228 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1016 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_988 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_966 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1006 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_207 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_229 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_218 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_390 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_978 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1018 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_208 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_219 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_391 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_380 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_968 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_209 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1008 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_392 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_370 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_381 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_371 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_393 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_360 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_382 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_190 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_394 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_350 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_372 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_361 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_383 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_191 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_180 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_395 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_351 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_362 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_340 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_384 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_373 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_192 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_181 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_170 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_330 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_341 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_396 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_352 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_374 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_363 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_385 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_193 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_182 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_160 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_171 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_512 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_397 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_353 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_320 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_375 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_386 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_364 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_342 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_331 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_194 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_183 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_161 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_172 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_150 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_354 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_310 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_343 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_321 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_332 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_398 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_376 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_387 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_365 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_184 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_195 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_162 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_173 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_140 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_151 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_333 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_300 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_399 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_344 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_311 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_377 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_388 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_366 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_322 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_355 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_196 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_185 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_163 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_174 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_130 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_141 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_152 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_90 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_334 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_301 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_345 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_389 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_378 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_367 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_323 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_312 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_356 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_120 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_197 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_186 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_164 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_175 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_131 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_142 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_153 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_91 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_80 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_335 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_302 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_379 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_346 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_368 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_324 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_313 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_357 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_198 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_187 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_165 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_176 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_132 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_143 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_121 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_110 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_154 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_92 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_70 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_81 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_303 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_347 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_336 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_369 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_325 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_314 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_358 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_188 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_199 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_166 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_177 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_144 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_111 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_100 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_133 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_122 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_155 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_93 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_60 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_82 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_71 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_304 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_348 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_326 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_337 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_315 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_359 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_167 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_189 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_178 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_112 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_134 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_123 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_156 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_145 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_101 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_50 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_94 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_61 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_72 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_83 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_305 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_327 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_349 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_338 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_316 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_168 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_179 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_124 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_135 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_157 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_113 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_146 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_102 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_40 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_51 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_95 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_62 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_73 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_84 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_328 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_306 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_339 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_317 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_114 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_103 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_125 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_169 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_158 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_136 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_147 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_41 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_52 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_30 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_96 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_63 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_74 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_85 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_329 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_307 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_318 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_115 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_137 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_159 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_148 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_104 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_126 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_42 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_53 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_20 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_31 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_64 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_75 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_86 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_97 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_319 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_308 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_116 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_138 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_127 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_149 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_105 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_43 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_10 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_54 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_21 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_32 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_65 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_87 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_98 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_76 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_309 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_139 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_106 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_128 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_117 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_470 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_44 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_11 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_55 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_22 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_33 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_99 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_88 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_66 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_77 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_118 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_129 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_107 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_471 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_460 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_290 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_45 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_12 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_34 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_23 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_56 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_67 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_78 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_89 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_108 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_119 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_472 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_461 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_450 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_280 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_291 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_46 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_13 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_35 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_24 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_57 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_68 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_79 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_109 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_451 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_440 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_462 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_473 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_292 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_281 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_270 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_14 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_47 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_36 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_25 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_58 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_69 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_452 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_430 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_463 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_441 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_474 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_260 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_282 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_293 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_271 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_15 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_48 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_37 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_26 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_59 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_464 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_475 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_453 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_420 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_431 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_442 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_4 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_261 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_283 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_250 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_294 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_272 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_49 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_38 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_27 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_16 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_476 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_454 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_421 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_465 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_410 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_443 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_432 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_5 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_262 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_284 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_251 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_295 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_240 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_273 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_39 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_17 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_28 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_477 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_455 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_422 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_411 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_466 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_433 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_444 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_400 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_6 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_230 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_296 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_263 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_285 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_252 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_241 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_274 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_18 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_29 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_3v256x8m81 m3_82_330# a_248_342# a_62_178# w_30_512#
+ a_430_96# a_110_96# a_192_298# VSUBS
X0 a_192_298# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_408_342# a_248_342# a_192_298# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_408_342# a_248_342# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_408_342# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt pmos_5p04310591302095_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4251p pd=2.155u as=0.7194p ps=4.15u w=1.635u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7194p pd=4.15u as=0.4251p ps=2.155u w=1.635u l=0.28u
.ends

.subckt nmos_5p04310591302098_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1664p pd=1.16u as=0.2816p ps=2.16u w=0.64u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.2816p pd=2.16u as=0.1664p ps=1.16u w=0.64u l=0.28u
.ends

.subckt pmos_5p04310591302097_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.2909p pd=5.485u as=2.1846p ps=10.81u w=4.965u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=2.1846p pd=10.81u as=1.2909p ps=5.485u w=4.965u l=0.28u
.ends

.subckt ypass_gate_3v256x8m81_0 bb db ypass d pcb m3_0_2091# pmos_5p0431059130201_3v256x8m81_2/D
+ m3_0_2831# a_64_1295# m3_0_3056# pmos_5p0431059130201_3v256x8m81_0/D m3_0_3781#
+ m3_0_1632# vss m3_0_3536# b m3_0_3291# m3_0_2331# m3_0_2581# vdd
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D a_64_1295#
+ a_64_1295# vss vss nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd b pmos_5p0431059130201_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 b pcb vdd bb pmos_5p0431059130201_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_2 pmos_5p0431059130201_3v256x8m81_2/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v256x8m81
Xnmos_5p0431059130200_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_2/D a_64_1295#
+ bb vss nmos_5p0431059130200_3v256x8m81
Xnmos_5p0431059130200_3v256x8m81_1 pmos_5p0431059130201_3v256x8m81_0/D a_64_1295#
+ b vss nmos_5p0431059130200_3v256x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
X1 bb pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X2 nmos_5p0431059130202_3v256x8m81_0/D a_64_1295# vdd vdd pfet_03v3 ad=0.1946p pd=1.255u as=0.38225p ps=2.49u w=0.695u l=0.28u
X3 vdd a_64_1295# nmos_5p0431059130202_3v256x8m81_0/D vdd pfet_03v3 ad=0.50735p pd=2.85u as=0.1946p ps=1.255u w=0.695u l=0.28u
X4 b pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X5 vdd pcb bb vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
.ends

.subckt nmos_5p04310591302096_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=1.0309p pd=4.485u as=1.7446p ps=8.81u w=3.965u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=1.7446p pd=8.81u as=1.0309p ps=4.485u w=3.965u l=0.28u
.ends

.subckt rdummy_3v256x4_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_62/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512# ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_3v256x8m81_62/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ pmos_5p04310591302097_3v256x8m81_0/D m3_15667_n5798# 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_43/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_43/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_7/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/m3_82_330# w_15880_n13729#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_63/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_63/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_10/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_44/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_44/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_8/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_30/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_30/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ m1_16100_n16182# 018SRAM_cell1_dummy_3v256x8m81_54/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_54/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/a_248_342# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_64/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_11/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_35/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_35/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_45/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_9/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_55/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_12/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_12/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_36/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_36/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_46/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_56/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_342# m3_15667_n5552#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_13/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_37/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_37/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_47/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_47/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_33/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_0/a_248_342#
+ ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D 018SRAM_cell1_dummy_R_3v256x8m81_33/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_57/m2_346_89#
+ m3_15667_n6510# 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_57/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89#
+ ypass_gate_3v256x8m81_0_0/vdd 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_14/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_38/m2_346_89#
+ m3_15667_n6288# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_38/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ a_n547_1214# 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_15/m3_82_330# m3_15698_n15942# 018SRAM_cell1_dummy_R_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_39/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_39/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_25/a_248_342#
+ m3_15667_n7247# 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_35/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_59/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_59/m2_134_89#
+ a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_16/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_16/a_248_342# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_26/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/a_248_342# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# m3_15645_n13711# 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_17/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_17/a_248_342# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_27/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_27/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_40/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_40/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_4/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_50/m2_134_89# pmos_5p04310591302097_3v256x8m81_0/S
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_60/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_60/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_18/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_18/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/m3_82_330# m3_15667_n6043#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_28/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_28/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_41/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_41/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_5/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_51/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_61/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_61/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_32/m2_346_89#
+ pmos_5p04310591302095_3v256x8m81_0/S 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_32/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_29/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_29/a_248_342#
+ m3_15667_n7002# 018SRAM_cell1_dummy_3v256x8m81_42/m2_346_89# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_42/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_6/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v256x8m81_6/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_39/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_52/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# a_16524_19394# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ ypass_gate_3v256x8m81_0_0/pcb 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_52/m2_134_89#
+ m3_15667_n6752#
X018SRAM_cell1_2x_3v256x8m81_7 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_19 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_5 018SRAM_cell1_dummy_R_3v256x8m81_5/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_5/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_10 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_21 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_54 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_54/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_54/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_43 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_43/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_43/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_32 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_32/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_32/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_25 018SRAM_cell1_dummy_R_3v256x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_25/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_14 018SRAM_cell1_dummy_R_3v256x8m81_14/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_14/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_8 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_6 018SRAM_cell1_dummy_R_3v256x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_6/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_22 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_55 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_55/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_44 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_44/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_44/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_33 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_33/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_26 018SRAM_cell1_dummy_R_3v256x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_26/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_15 018SRAM_cell1_dummy_R_3v256x8m81_15/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_15/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
Xpmos_5p04310591302095_3v256x8m81_0 pmos_5p04310591302095_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/S
+ pmos_5p04310591302095_3v256x8m81_0/S pmos_5p04310591302095_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_7 018SRAM_cell1_dummy_R_3v256x8m81_7/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_7/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_23 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_56 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_56/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_45 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_45/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_34 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_34/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_38 018SRAM_cell1_dummy_R_3v256x8m81_38/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_27 018SRAM_cell1_dummy_R_3v256x8m81_27/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_27/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_16 018SRAM_cell1_dummy_R_3v256x8m81_16/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_16/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_8 018SRAM_cell1_dummy_R_3v256x8m81_8/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_8/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_24 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_57 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_57/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_57/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_46 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_46/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_35 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_35/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_35/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_39 018SRAM_cell1_dummy_R_3v256x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_39/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_28 018SRAM_cell1_dummy_R_3v256x8m81_28/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_28/a_248_342# a_16524_19394# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_17 018SRAM_cell1_dummy_R_3v256x8m81_17/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_17/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_9 018SRAM_cell1_dummy_R_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_9/a_248_342# a_16524_2# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_25 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_47 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_47/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_47/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_36 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_36/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_36/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_29 018SRAM_cell1_dummy_R_3v256x8m81_29/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_29/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_18 018SRAM_cell1_dummy_R_3v256x8m81_18/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_18/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_26 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_59 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_59/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_59/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_48 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_48/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_37 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_37/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_37/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_19 a_n547_48# ypass_gate_3v256x8m81_0_0/vss a_16524_2#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_16 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_27 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_49 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_49/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_38 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_38/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_38/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_17 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_28 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_39 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_39/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_39/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
Xnmos_5p04310591302098_3v256x8m81_0 pmos_5p04310591302095_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/vss
+ ypass_gate_3v256x8m81_0_0/vss nmos_5p04310591302098_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_18 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_29 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_19 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_0 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ a_n547_48# 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
Xpmos_5p04310591302097_3v256x8m81_0 pmos_5p04310591302097_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/D
+ pmos_5p04310591302095_3v256x8m81_0/D w_15880_n13729# pmos_5p04310591302097_3v256x8m81_0/S
+ pmos_5p04310591302097_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ a_n547_1214# 018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
Xypass_gate_3v256x8m81_0_0 ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/db
+ ypass_gate_3v256x8m81_0_0/ypass ypass_gate_3v256x8m81_0_0/d ypass_gate_3v256x8m81_0_0/pcb
+ m3_15667_n7247# ypass_gate_3v256x8m81_0_0/bb m3_15667_n6510# ypass_gate_3v256x8m81_0_0/vdd
+ m3_15667_n6288# ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D m3_15667_n5552#
+ ypass_gate_3v256x8m81_0_0/vdd ypass_gate_3v256x8m81_0_0/vss m3_15667_n5798# ypass_gate_3v256x8m81_0_0/b
+ m3_15667_n6043# m3_15667_n7002# m3_15667_n6752# ypass_gate_3v256x8m81_0_0/vdd ypass_gate_3v256x8m81_0
X018SRAM_cell1_dummy_3v256x8m81_4 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_31 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
Xnmos_5p04310591302096_3v256x8m81_0 pmos_5p04310591302097_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/D
+ pmos_5p04310591302095_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/vss ypass_gate_3v256x8m81_0_0/vss
+ nmos_5p04310591302096_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_40 018SRAM_cell1_dummy_R_3v256x8m81_40/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_52 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss
+ a_16524_19394# 018SRAM_cell1_3v256x8m81_1/w_30_512# ypass_gate_3v256x8m81_0_0/bb
+ ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_1/w_30_512# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_30 018SRAM_cell1_dummy_R_3v256x8m81_30/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_30/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_0 018SRAM_cell1_dummy_R_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_14 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_60 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_60/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_60/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_1 018SRAM_cell1_dummy_R_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_15 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_61 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_61/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_61/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_50 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_50/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_65 018SRAM_cell1_dummy_R_3v256x8m81_65/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_10 018SRAM_cell1_dummy_R_3v256x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_10/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_4 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_2 018SRAM_cell1_dummy_R_3v256x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_16 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_62 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_62/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_62/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_51 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_51/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_40 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_40/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_40/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_33 018SRAM_cell1_dummy_R_3v256x8m81_33/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_33/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_11 018SRAM_cell1_dummy_R_3v256x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_11/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_5 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_3 018SRAM_cell1_dummy_R_3v256x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_17 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_30 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_63 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_63/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_63/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_52 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_52/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_52/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_41 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_41/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_41/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_34 018SRAM_cell1_dummy_R_3v256x8m81_34/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_12 018SRAM_cell1_dummy_R_3v256x8m81_12/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_12/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_6 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_4 018SRAM_cell1_dummy_R_3v256x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_18 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# a_n547_1214# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# a_n547_1214# ypass_gate_3v256x8m81_0_0/vss
+ x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_20 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_31 a_n547_48# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_48# 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_64 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_64/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_53 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_53/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_42 a_16524_19394# ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# a_16524_19394# 018SRAM_cell1_dummy_3v256x8m81_42/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_42/m2_134_89# ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_35 018SRAM_cell1_dummy_R_3v256x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_35/a_248_342# a_16524_19394# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_13 018SRAM_cell1_dummy_R_3v256x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_13/a_248_342# a_16524_2# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ ypass_gate_3v256x8m81_0_0/vss x018SRAM_cell1_dummy_R_3v256x8m81
.ends

.subckt rcol4_256_3v256x8m81 WL[29] WL[20] WL[27] WL[30] WL[18] WL[15] WL[31] WL[14]
+ WL[16] WL[26] WL[19] WL[28] WL[12] WL[8] WL[5] WL[10] WL[13] WL[6] tblhl GWE WL[11]
+ din[7] q[5] q[6] q[7] din[5] din[6] q[4] pcb[7] pcb[4] WEN[4] WEN[7] pcb[5] WEN[5]
+ WEN[6] rarray4_256_3v256x8m81_0/m3_n1397_10705# rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/pcb
+ rarray4_256_3v256x8m81_0/m3_n1397_8779# rarray4_256_3v256x8m81_0/m3_n1397_8281#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass saout_m2_3v256x8m81_3/din_3v256x8m81_0/men
+ saout_R_m2_3v256x8m81_1/datain saout_m2_3v256x8m81_2/q rarray4_256_3v256x8m81_0/m3_n1397_13129#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass rarray4_256_3v256x8m81_0/m3_n1397_11917#
+ rarray4_256_3v256x8m81_0/m3_n1397_9493# saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ rarray4_256_3v256x8m81_0/m3_n1397_5143# WL[21] WL[7] rarray4_256_3v256x8m81_0/m3_n1397_3931#
+ WL[1] WL[0] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ rarray4_256_3v256x8m81_0/m3_n1397_19687# rarray4_256_3v256x8m81_0/m3_n1397_6355#
+ WL[9] WL[23] WL[22] saout_m2_3v256x8m81_3/ypass[7] saout_R_m2_3v256x8m81_1/q saout_m2_3v256x8m81_3/q
+ WL[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass rdummy_3v256x4_3v256x8m81_0/a_16524_2#
+ saout_R_m2_3v256x8m81_3/q saout_R_m2_3v256x8m81_3/datain rarray4_256_3v256x8m81_0/m3_n1397_7567#
+ WL[25] saout_m2_3v256x8m81_3/GWEN saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ WL[24] WL[4] WL[3] WL[17] pcb[6] VSS
Xrarray4_256_3v256x8m81_0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[17] saout_m2_3v256x8m81_3/bb[3] rarray4_256_3v256x8m81_0/m3_n1397_13129# saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_2/bb[5] WL[4] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ rarray4_256_3v256x8m81_0/m3_n1397_11917# saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_2/b[4] saout_R_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/b[4]
+ rarray4_256_3v256x8m81_0/m3_n1397_8779# saout_m2_3v256x8m81_2/bb[3] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[28] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_m2_3v256x8m81_3/b[3]
+ saout_R_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_1/b[3] WL[26] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ rarray4_256_3v256x8m81_0/m3_n1397_3931# WL[5] saout_R_m2_3v256x8m81_1/b[6] WL[3]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb WL[1] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ rarray4_256_3v256x8m81_0/m3_n1397_8281# saout_R_m2_3v256x8m81_1/bb[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[30] rarray4_256_3v256x8m81_0/m3_n1397_19687# saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/b[3]
+ WL[29] WL[15] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_2/b[3] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_3/bb[4] saout_m2_3v256x8m81_3/bb[2] WL[19] WL[23] WL[24] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb rarray4_256_3v256x8m81_0/m3_n1397_10705#
+ saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb WL[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_3/bb[7] WL[21] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[0] WL[2] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_1/bb[5]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_2/b[1]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_R_m2_3v256x8m81_1/bb[2] rarray4_256_3v256x8m81_0/m3_n1397_5143# rarray4_256_3v256x8m81_0/m3_n1397_9493#
+ WL[27] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/b[6]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[22] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb rarray4_256_3v256x8m81_0/m3_n1397_6355#
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_2/b[6] saout_R_m2_3v256x8m81_1/bb[4] rarray4_256_3v256x8m81_0/m3_n1397_7567#
+ pcb[6] WL[25] WL[11] saout_m2_3v256x8m81_2/bb[2] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ WL[9] VSS rarray4_256_3v256x8m81
Xrdummy_3v256x4_3v256x8m81_0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb pcb[6] rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b pcb[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[30] VSS tblhl saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ pcb[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b pcb[6]
+ saout_m2_3v256x8m81_3/bb[5] pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_7567# VSS saout_R_m2_3v256x8m81_3/bb[4]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b rarray4_256_3v256x8m81_0/m3_n1397_8779#
+ VSS saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_8779# pcb[6] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b saout_R_m2_3v256x8m81_1/bb[7]
+ VSS saout_m2_3v256x8m81_2/b[4] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[1] pcb[6] saout_R_m2_3v256x8m81_1/bb[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ WL[5] VSS pcb[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[25] pcb[6] VSS saout_m2_3v256x8m81_3/b[4] pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_8281#
+ VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/bb[5]
+ rarray4_256_3v256x8m81_0/m3_n1397_7567# WL[25] VSS VSS pcb[6] pcb[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ rarray4_256_3v256x8m81_0/m3_n1397_9493# tblhl saout_m2_3v256x8m81_2/b[3] saout_R_m2_3v256x8m81_1/b[6]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb VSS saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_2/bb[3] WL[28] WL[17] VSS VSS pcb[6] saout_R_m2_3v256x8m81_1/bb[2]
+ saout_m2_3v256x8m81_3/bb[2] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b WL[7] pcb[6]
+ VSS pcb[6] pcb[6] WL[26] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSS saout_m2_3v256x8m81_3/b[6] pcb[6] saout_R_m2_3v256x8m81_3/b[3] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[0] VSS pcb[6] pcb[6] saout_m2_3v256x8m81_2/bb[2] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/b[6]
+ rarray4_256_3v256x8m81_0/m3_n1397_6355# rarray4_256_3v256x8m81_0/m3_n1397_11917#
+ VSS VSS saout_m2_3v256x8m81_3/b[3] saout_m2_3v256x8m81_3/bb[3] WL[11] pcb[6] VSS
+ pcb[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ pcb[6] pcb[6] WL[23] VSS saout_R_m2_3v256x8m81_3/bb[2] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ pcb[6] pcb[6] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/bb[4]
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ WL[11] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b pcb[6] pcb[6]
+ saout_m2_3v256x8m81_3/bb[5] pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_9493# VSS pcb[6]
+ saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ pcb[6] WL[24] VSS pcb[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_3931# WL[22] VSS rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/b
+ VSS saout_m2_3v256x8m81_2/b[1] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb saout_R_m2_3v256x8m81_3/bb[5]
+ saout_R_m2_3v256x8m81_1/b[6] pcb[6] WL[15] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VSS pcb[6] saout_m2_3v256x8m81_3/b[4] pcb[6] pcb[6] WL[3] VSS pcb[6] saout_m2_3v256x8m81_3/bb[2]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass WL[0] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b WL[27] saout_m2_3v256x8m81_2/bb[5]
+ VSS rarray4_256_3v256x8m81_0/m3_n1397_5143# pcb[6] WL[26] VSS VSS saout_m2_3v256x8m81_2/bb[2]
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/b[3]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb rarray4_256_3v256x8m81_0/m3_n1397_10705#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb VSS VSS pcb[6]
+ saout_m2_3v256x8m81_3/b[6] WL[9] VSS VSS pcb[6] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ WL[1] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb VSS
+ WL[23] pcb[6] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ pcb[6] pcb[6] saout_m2_3v256x8m81_2/b[1] WL[28] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VSS WL[4] WL[30] VSS VSS saout_m2_3v256x8m81_2/b[3] pcb[6] saout_R_m2_3v256x8m81_1/b[3]
+ saout_m2_3v256x8m81_2/bb[3] pcb[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ rdummy_3v256x4_3v256x8m81_0/a_16524_2# rarray4_256_3v256x8m81_0/m3_n1397_8281# rarray4_256_3v256x8m81_0/m3_n1397_5143#
+ VSS VSS rarray4_256_3v256x8m81_0/m3_n1397_11917# WL[19] VSS VSS pcb[6] rarray4_256_3v256x8m81_0/m3_n1397_3931#
+ VSS WL[2] VSS WL[19] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ pcb[6] pcb[6] VSS saout_R_m2_3v256x8m81_1/bb[4] saout_m2_3v256x8m81_2/bb[5] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ WL[21] saout_R_m2_3v256x8m81_3/bb[2] VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ rarray4_256_3v256x8m81_0/m3_n1397_10705# WL[9] VSS VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb WL[21] VSS
+ pcb[6] WL[7] VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/bb[7] rarray4_256_3v256x8m81_0/m3_n1397_6355# pcb[6] VSS
+ rarray4_256_3v256x8m81_0/m3_n1397_13129# saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b pcb[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_2/b[4] saout_R_m2_3v256x8m81_1/bb[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ pcb[6] pcb[6] WL[22] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b VSS pcb[6]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ WL[1] pcb[6] VSS pcb[6] pcb[6] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[4] saout_m2_3v256x8m81_3/ypass[7] VSS saout_R_m2_3v256x8m81_3/bb[7] WL[29] VSS
+ pcb[6] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[2] VSS WL[17] rarray4_256_3v256x8m81_0/m3_n1397_13129# VSS VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/b[3] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_2/b[6] pcb[6] saout_m2_3v256x8m81_2/b[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VSS saout_R_m2_3v256x8m81_1/bb[4] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[29] VSS pcb[6] saout_m2_3v256x8m81_3/b[3] pcb[6] WL[5] saout_m2_3v256x8m81_3/bb[3]
+ VSS WL[27] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb pcb[6] saout_R_m2_3v256x8m81_3/b[6]
+ WL[3] VSS WL[24] WL[15] pcb[6] VSS VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ VSS pcb[6] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_R_m2_3v256x8m81_1/bb[2] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ rarray4_256_3v256x8m81_0/m3_n1397_19687# pcb[6] rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/pcb
+ pcb[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass rdummy_3v256x4_3v256x8m81
Xsaout_R_m2_3v256x8m81_1 saout_R_m2_3v256x8m81_1/ypass[2] saout_R_m2_3v256x8m81_1/ypass[3]
+ saout_R_m2_3v256x8m81_1/ypass[4] saout_R_m2_3v256x8m81_1/ypass[5] saout_R_m2_3v256x8m81_1/ypass[6]
+ GWE saout_m2_3v256x8m81_3/GWEN saout_R_m2_3v256x8m81_1/datain saout_R_m2_3v256x8m81_1/b[5]
+ saout_R_m2_3v256x8m81_1/b[4] saout_R_m2_3v256x8m81_1/b[2] saout_R_m2_3v256x8m81_1/b[1]
+ saout_R_m2_3v256x8m81_1/b[0] saout_R_m2_3v256x8m81_1/bb[6] saout_R_m2_3v256x8m81_1/q
+ saout_R_m2_3v256x8m81_1/bb[3] saout_R_m2_3v256x8m81_1/bb[0] saout_R_m2_3v256x8m81_1/bb[1]
+ saout_R_m2_3v256x8m81_1/pcb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb WEN[4]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_1/bb[2]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/b[3]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass saout_m2_3v256x8m81_3/din_3v256x8m81_0/men
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_R_m2_3v256x8m81_1/bb[4]
+ saout_R_m2_3v256x8m81_1/b[6] saout_m2_3v256x8m81_3/ypass[7] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass saout_R_m2_3v256x8m81_1/bb[7]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ VSS pcb[6] saout_R_m2_3v256x8m81
Xsaout_R_m2_3v256x8m81_3 saout_R_m2_3v256x8m81_3/ypass[2] saout_R_m2_3v256x8m81_3/ypass[3]
+ saout_R_m2_3v256x8m81_3/ypass[4] saout_R_m2_3v256x8m81_3/ypass[5] saout_R_m2_3v256x8m81_3/ypass[6]
+ GWE saout_m2_3v256x8m81_3/GWEN saout_R_m2_3v256x8m81_3/datain saout_R_m2_3v256x8m81_3/b[5]
+ saout_R_m2_3v256x8m81_3/b[4] saout_R_m2_3v256x8m81_3/b[2] saout_R_m2_3v256x8m81_3/b[1]
+ saout_R_m2_3v256x8m81_3/b[0] saout_R_m2_3v256x8m81_3/bb[6] saout_R_m2_3v256x8m81_3/q
+ saout_R_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_3/bb[0] saout_R_m2_3v256x8m81_3/bb[1]
+ saout_R_m2_3v256x8m81_3/pcb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/sa_3v256x8m81_0/pcb WEN[6]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_3/bb[2]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_3/b[3]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass saout_m2_3v256x8m81_3/din_3v256x8m81_0/men
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_R_m2_3v256x8m81_3/bb[4]
+ saout_R_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/ypass[7] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass saout_R_m2_3v256x8m81_3/bb[7]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ VSS pcb[6] saout_R_m2_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[0] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[1] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[2] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[3] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[4] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[5] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[6] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[7] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[8] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[9] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[10] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[11] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[12] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[13] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[14] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[15] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[16] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[17] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[18] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[19] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[20] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[21] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[22] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[23] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[24] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[25] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[26] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[27] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[28] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[29] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[30] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[31] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[32] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[33] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[34] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[35] pcb[6] VSS pcb[6] dcap_103_novia_3v256x8m81
Xsaout_m2_3v256x8m81_2 saout_m2_3v256x8m81_2/ypass[2] saout_m2_3v256x8m81_2/ypass[3]
+ saout_m2_3v256x8m81_2/ypass[4] saout_m2_3v256x8m81_2/ypass[5] saout_m2_3v256x8m81_2/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN GWE saout_m2_3v256x8m81_2/bb[1] saout_m2_3v256x8m81_2/bb[4]
+ saout_m2_3v256x8m81_2/bb[7] saout_m2_3v256x8m81_2/bb[6] saout_m2_3v256x8m81_2/b[5]
+ saout_m2_3v256x8m81_2/b[7] saout_m2_3v256x8m81_2/b[2] saout_m2_3v256x8m81_2/q saout_m2_3v256x8m81_2/pcb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_2/b[6] saout_m2_3v256x8m81_2/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ WEN[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/bb[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_2/b[4] saout_m2_3v256x8m81_3/din_3v256x8m81_0/men saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ GWE saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_2/bb[3] saout_m2_3v256x8m81_2/b[1] saout_m2_3v256x8m81_3/ypass[7]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass saout_m2_3v256x8m81_2/b[3]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ pcb[6] saout_m2_3v256x8m81
Xsaout_m2_3v256x8m81_3 saout_m2_3v256x8m81_3/ypass[2] saout_m2_3v256x8m81_3/ypass[3]
+ saout_m2_3v256x8m81_3/ypass[4] saout_m2_3v256x8m81_3/ypass[5] saout_m2_3v256x8m81_3/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN GWE saout_m2_3v256x8m81_3/bb[1] saout_m2_3v256x8m81_3/bb[4]
+ saout_m2_3v256x8m81_3/bb[7] saout_m2_3v256x8m81_3/bb[6] saout_m2_3v256x8m81_3/b[5]
+ saout_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[2] saout_m2_3v256x8m81_3/q saout_m2_3v256x8m81_3/pcb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ WEN[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_3/bb[5] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_3/b[4] saout_m2_3v256x8m81_3/din_3v256x8m81_0/men saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ GWE saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_3/bb[3] saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/ypass[7]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass saout_m2_3v256x8m81_3/b[3]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ pcb[6] saout_m2_3v256x8m81
.ends

.subckt pmos_5p04310591302058_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.9306p pd=5.11u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$47331372_3v256x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302058_3v256x8m81_0/S
+ a_118_n34# pmos_5p04310591302058_3v256x8m81_0/D
Xpmos_5p04310591302058_3v256x8m81_0 pmos_5p04310591302058_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302058_3v256x8m81_0/S pmos_5p04310591302058_3v256x8m81
.ends

.subckt pmos_1p2_160_3v256x8m81 w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81_0/D
+ a_n14_n34#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt nmos_5p04310591302059_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.28u
.ends

.subckt nmos_1p2$$47329324_3v256x8m81 a_118_n34# a_n41_n34# nmos_5p04310591302059_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302059_3v256x8m81_0/D
Xnmos_5p04310591302059_3v256x8m81_0 nmos_5p04310591302059_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302059_3v256x8m81_0/S VSUBS nmos_5p04310591302059_3v256x8m81
.ends

.subckt pmos_1p2_161_3v256x8m81 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89# pmos_5p04310591302041_3v256x8m81_0/S
+ w_n133_n65#
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
.ends

.subckt nmos_1p2_157_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34# nmos_5p04310591302010_3v256x8m81_0/S
+ VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt alatch_3v256x8m81 enb en ab a a_886_665# vdd vss
Xpmos_1p2$$47331372_3v256x8m81_0 pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ vdd vdd pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S ab pmos_1p2$$47331372_3v256x8m81
Xpmos_1p2_160_3v256x8m81_0 vdd pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ a enb pmos_1p2_160_3v256x8m81
Xnmos_1p2$$47329324_3v256x8m81_0 pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S vss vss ab nmos_1p2$$47329324_3v256x8m81
Xpmos_1p2_161_3v256x8m81_0 pmos_1p2_161_3v256x8m81_1/pmos_5p04310591302041_3v256x8m81_0/S
+ a_886_665# pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S vdd pmos_1p2_161_3v256x8m81
Xpmos_1p2_161_3v256x8m81_1 vdd ab pmos_1p2_161_3v256x8m81_1/pmos_5p04310591302041_3v256x8m81_0/S
+ vdd pmos_1p2_161_3v256x8m81
Xnmos_1p2_157_3v256x8m81_0 a a_886_665# pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ vss nmos_1p2_157_3v256x8m81
X0 pmos_1p2_161_3v256x8m81_1/pmos_5p04310591302041_3v256x8m81_0/S enb pmos_1p2_161_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss ab pmos_1p2_161_3v256x8m81_1/pmos_5p04310591302041_3v256x8m81_0/S vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302057_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.9306p pd=5.11u as=0.9306p ps=5.11u w=2.115u l=0.28u
.ends

.subckt nmos_1p2$$47514668_3v256x8m81 nmos_5p04310591302057_3v256x8m81_0/S nmos_5p04310591302057_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v256x8m81_0 nmos_5p04310591302057_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v256x8m81_0/S VSUBS nmos_5p04310591302057_3v256x8m81
.ends

.subckt ypredec1_bot_3v256x8m81 m1_n9_2295# m1_n9_2436# m1_n9_2154# alatch_3v256x8m81_0/a
+ m1_n9_2013# m1_n9_1871# pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ m1_n9_1730# pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/enb alatch_3v256x8m81_0/vss pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ m2_800_896#
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/enb alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab
+ alatch_3v256x8m81_0/a m2_800_896# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/vss
+ alatch_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_0 alatch_3v256x8m81_0/vss pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D alatch_3v256x8m81_0/vss
+ nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_1 alatch_3v256x8m81_0/vss pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ alatch_3v256x8m81_0/ab alatch_3v256x8m81_0/vss nmos_1p2$$47514668_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_0 pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D pmos_1p2$$46887980_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_1 pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S alatch_3v256x8m81_0/ab
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D pmos_1p2$$46887980_3v256x8m81
.ends

.subckt pmos_5p04310591302055_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.1052p pd=19.54u as=4.1052p ps=19.54u w=9.33u l=0.28u
.ends

.subckt nmos_5p04310591302054_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.8634p pd=9.35u as=1.8634p ps=9.35u w=4.235u l=0.28u
.ends

.subckt ypredec1_ys_3v256x8m81 a_161_1551# nmos_5p04310591302054_3v256x8m81_1/D pmos_5p04310591302055_3v256x8m81_1/S
+ pmos_5p04310591302055_3v256x8m81_3/S nmos_5p04310591302054_3v256x8m81_2/S nmos_5p04310591302054_3v256x8m81_3/D
+ pmos_5p04310591302055_3v256x8m81_3/D VSUBS
Xpmos_5p04310591302055_3v256x8m81_0 pmos_5p04310591302055_3v256x8m81_0/D a_161_1551#
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_1 pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_1/S pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_2 pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_3 pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_0 pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81_0/D
+ nmos_5p04310591302054_3v256x8m81_1/D VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_1 nmos_5p04310591302054_3v256x8m81_1/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_1/S VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_2 pmos_5p04310591302055_3v256x8m81_0/D a_161_1551#
+ nmos_5p04310591302054_3v256x8m81_2/S VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_3 nmos_5p04310591302054_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/S VSUBS nmos_5p04310591302054_3v256x8m81
.ends

.subckt nmos_5p04310591302056_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3916p pd=2.66u as=0.3916p ps=2.66u w=0.89u l=0.28u
.ends

.subckt nmos_1p2$$47342636_3v256x8m81 a_n14_n44# a_n102_0# a_42_0# VSUBS
X0 a_42_0# a_n14_n44# a_n102_0# VSUBS nfet_03v3 ad=0.2772p pd=2.14u as=0.2772p ps=2.14u w=0.63u l=0.28u
.ends

.subckt pmos_5p04310591302061_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1836p pd=6.26u as=1.1836p ps=6.26u w=2.69u l=0.28u
.ends

.subckt pmos_1p2$$47820844_3v256x8m81 pmos_5p04310591302061_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302061_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302061_3v256x8m81_0 pmos_5p04310591302061_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302061_3v256x8m81_0/S pmos_5p04310591302061_3v256x8m81
.ends

.subckt pmos_5p04310591302060_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1638p pd=6.17u as=1.1638p ps=6.17u w=2.645u l=0.28u
.ends

.subckt pmos_1p2$$47821868_3v256x8m81 pmos_5p04310591302060_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302060_3v256x8m81_0/D w_n133_n66#
Xpmos_5p04310591302060_3v256x8m81_0 pmos_5p04310591302060_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302060_3v256x8m81_0/S pmos_5p04310591302060_3v256x8m81
.ends

.subckt ypredec1_xa_3v256x8m81 m1_n40_n2861# a_145_n4683# m3_0_n4986# m1_n40_n3567#
+ m1_n40_n3285# pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# a_0_56# a_465_n4683# m1_n40_n3426#
+ m1_n40_n3144# pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# M2_M1$$47515692_3v256x8m81_0/VSUBS
+ pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D m1_n40_n3003#
+ a_305_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
Xpmos_1p2$$47820844_3v256x8m81_0 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47820844_3v256x8m81_1 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47820844_3v256x8m81_2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_0 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ a_145_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 M2_M1$$47515692_3v256x8m81_0/VSUBS pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D M2_M1$$47515692_3v256x8m81_0/VSUBS
+ nmos_1p2$$46551084_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_1 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D M2_M1$$47515692_3v256x8m81_0/VSUBS
+ M2_M1$$47515692_3v256x8m81_0/VSUBS nmos_1p2$$46551084_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ a_305_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_2 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D M2_M1$$47515692_3v256x8m81_0/VSUBS
+ M2_M1$$47515692_3v256x8m81_0/VSUBS nmos_1p2$$46551084_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_3 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ a_465_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
X0 a_361_n4624# a_305_n4683# a_201_n4624# M2_M1$$47515692_3v256x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=0.8268p ps=3.7u w=3.18u l=0.28u
X1 a_201_n4624# a_145_n4683# M2_M1$$47515692_3v256x8m81_0/VSUBS M2_M1$$47515692_3v256x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=1.4469p ps=7.27u w=3.18u l=0.28u
X2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D a_465_n4683# a_361_n4624# M2_M1$$47515692_3v256x8m81_0/VSUBS nfet_03v3 ad=1.5423p pd=7.33u as=0.8268p ps=3.7u w=3.18u l=0.28u
.ends

.subckt ypredec1_xax8_3v256x8m81 ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_997_2070# ypredec1_xa_3v256x8m81_3/a_0_56# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_683_1364# ypredec1_xa_3v256x8m81_5/a_0_56# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ a_4427_1646# ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_4270_1505# VSUBS a_526_1788#
Xypredec1_xa_3v256x8m81_0 a_997_2070# a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_0/a_0_56# a_4427_1646# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_840_1930# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_1 a_997_2070# a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_5/a_0_56# a_4427_1646# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_4270_1505# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_2 a_997_2070# a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ VSUBS a_997_2070# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_4270_1505# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_3 a_997_2070# a_526_1788# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_3/a_0_56# a_997_2070# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_840_1930# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_4 a_997_2070# a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_4/a_0_56# a_4427_1646# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_840_1930# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_5 a_997_2070# a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_5/a_0_56# a_4427_1646# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_4270_1505# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_6 a_997_2070# a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_6/a_0_56# a_997_2070# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_4270_1505# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_7 a_997_2070# a_683_1364# VSUBS a_683_1364# a_4427_1646# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65#
+ ypredec1_xa_3v256x8m81_7/a_0_56# a_997_2070# a_4270_1505# a_526_1788# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ a_840_1930# a_840_1930# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
.ends

.subckt pmos_5p04310591302062_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$47109164_3v256x8m81 pmos_5p04310591302062_3v256x8m81_0/D pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ a_118_159# pmos_5p04310591302062_3v256x8m81_0/S a_n42_159#
Xpmos_5p04310591302062_3v256x8m81_0 pmos_5p04310591302062_3v256x8m81_0/D a_n42_159#
+ a_118_159# pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# pmos_5p04310591302062_3v256x8m81_0/S
+ pmos_5p04310591302062_3v256x8m81
.ends

.subckt ypredec1_3v256x8m81 ly[5] ly[4] ly[7] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/a
+ ly[3] ypredec1_bot_3v256x8m81_0/alatch_3v256x8m81_0/a pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ ypredec1_bot_3v256x8m81_1/alatch_3v256x8m81_0/a pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
Xypredec1_bot_3v256x8m81_1 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_4 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[0] ly[0] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_bot_3v256x8m81_2 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_5 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[1] ly[1] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_6 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[2] ly[2] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_7 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[5] ry[5] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_8 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[6] ry[6] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_9 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[7] ry[7] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_10 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[1] ry[1] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_11 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[2] ry[2] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_12 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[3] ry[3] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_0 M1_NWELL13_3v256x8m81_0/VSUBS clk nmos_5p04310591302056_3v256x8m81_1/D
+ M1_NWELL13_3v256x8m81_0/VSUBS nmos_5p04310591302056_3v256x8m81
Xypredec1_ys_3v256x8m81_13 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[4] ry[4] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_1 nmos_5p04310591302056_3v256x8m81_1/D men M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS nmos_5p04310591302056_3v256x8m81
Xypredec1_ys_3v256x8m81_14 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[0] ry[0] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_15 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[7] ly[7] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS nmos_1p2$$47342636_3v256x8m81
Xypredec1_xax8_3v256x8m81_0 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81
Xypredec1_ys_3v256x8m81_0 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[3] ly[3] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_1 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[4] ly[4] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xpmos_1p2$$47109164_3v256x8m81_0 ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# nmos_5p04310591302056_3v256x8m81_1/D
+ pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S nmos_5p04310591302056_3v256x8m81_1/D
+ pmos_1p2$$47109164_3v256x8m81
Xypredec1_ys_3v256x8m81_2 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[5] ly[5] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_bot_3v256x8m81_0 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_3 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[6] ly[6] M1_NWELL13_3v256x8m81_0/VSUBS M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
X0 a_5490_186# clk nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.1917p pd=1.425u as=0.34345p ps=1.71u w=1.065u l=0.28u
X1 nmos_5p04310591302056_3v256x8m81_1/D clk a_5176_186# pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.34345p pd=1.71u as=0.19435p ps=1.43u w=1.065u l=0.28u
X2 a_5176_186# men pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.19435p pd=1.43u as=0.59108p ps=3.24u w=1.065u l=0.28u
X3 pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S men a_5490_186# pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.59108p pd=3.24u as=0.1917p ps=1.425u w=1.065u l=0.28u
.ends

.subckt pmos_5p04310591302068_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt pmos_1p2$$47513644_3v256x8m81 pmos_5p04310591302068_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302068_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302068_3v256x8m81_0 pmos_5p04310591302068_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302068_3v256x8m81_0/S pmos_5p04310591302068_3v256x8m81
.ends

.subckt pmos_5p04310591302072_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.1406p pd=10.61u as=2.1406p ps=10.61u w=4.865u l=0.28u
.ends

.subckt pmos_1p2$$47512620_3v256x8m81 a_n14_n34# pmos_5p04310591302072_3v256x8m81_0/S
+ w_n133_n66# pmos_5p04310591302072_3v256x8m81_0/D
Xpmos_5p04310591302072_3v256x8m81_0 pmos_5p04310591302072_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302072_3v256x8m81_0/S pmos_5p04310591302072_3v256x8m81
.ends

.subckt xpredec1_xa_3v256x8m81 m1_n40_n4147# m1_n40_n4005# m3_n46_n5510# a_145_n5643#
+ m1_n40_n3864# m1_n40_n3582# m1_n40_n3723# a_0_56# m1_n40_n3441# a_465_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ M2_M1$$47515692_3v256x8m81_3/VSUBS a_305_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
Xpmos_1p2$$47513644_3v256x8m81_0 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_0 M2_M1$$47515692_3v256x8m81_3/VSUBS pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S M2_M1$$47515692_3v256x8m81_3/VSUBS
+ nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ M2_M1$$47515692_3v256x8m81_3/VSUBS pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ M2_M1$$47515692_3v256x8m81_3/VSUBS nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_2 M2_M1$$47515692_3v256x8m81_3/VSUBS pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S M2_M1$$47515692_3v256x8m81_3/VSUBS
+ nmos_1p2$$47514668_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_0 a_145_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_1 a_465_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_3 a_305_n5643# pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
X0 a_361_n5592# a_305_n5643# a_201_n5592# M2_M1$$47515692_3v256x8m81_3/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=1.5145p ps=6.345u w=5.825u l=0.28u
X1 a_201_n5592# a_145_n5643# M2_M1$$47515692_3v256x8m81_3/VSUBS M2_M1$$47515692_3v256x8m81_3/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=2.65037p ps=12.56u w=5.825u l=0.28u
X2 pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S a_465_n5643# a_361_n5592# M2_M1$$47515692_3v256x8m81_3/VSUBS nfet_03v3 ad=2.82512p pd=12.62u as=1.5145p ps=6.345u w=5.825u l=0.28u
.ends

.subckt nmos_5p04310591302071_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.3508p pd=7.02u as=1.3508p ps=7.02u w=3.07u l=0.28u
.ends

.subckt nmos_1p2$$47336492_3v256x8m81 nmos_5p04310591302071_3v256x8m81_0/S nmos_5p04310591302071_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302071_3v256x8m81_0 nmos_5p04310591302071_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302071_3v256x8m81_0/S VSUBS nmos_5p04310591302071_3v256x8m81
.ends

.subckt pmos_5p04310591302070_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.3528p pd=16.12u as=3.3528p ps=16.12u w=7.62u l=0.28u
.ends

.subckt pmos_1p2$$47337516_3v256x8m81 pmos_5p04310591302070_3v256x8m81_0/S pmos_5p04310591302070_3v256x8m81_0/D
+ a_n14_n34# w_n133_n65#
Xpmos_5p04310591302070_3v256x8m81_0 pmos_5p04310591302070_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302070_3v256x8m81_0/S pmos_5p04310591302070_3v256x8m81
.ends

.subckt xpredec1_bot_3v256x8m81 m1_n74_2740# pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ alatch_3v256x8m81_0/a pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ m1_n74_3446# alatch_3v256x8m81_0/enb m1_n74_3164# m2_800_1786# m1_n74_3305# m1_n74_3023#
+ alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/vss pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ m1_n74_2881#
Xnmos_1p2$$47336492_3v256x8m81_0 alatch_3v256x8m81_0/vss pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D alatch_3v256x8m81_0/vss
+ nmos_1p2$$47336492_3v256x8m81
Xnmos_1p2$$47336492_3v256x8m81_1 alatch_3v256x8m81_0/vss pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ alatch_3v256x8m81_0/ab alatch_3v256x8m81_0/vss nmos_1p2$$47336492_3v256x8m81
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/enb alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab
+ alatch_3v256x8m81_0/a m2_800_1786# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/vss
+ alatch_3v256x8m81
Xpmos_1p2$$47337516_3v256x8m81_0 pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S pmos_1p2$$47337516_3v256x8m81
Xpmos_1p2$$47337516_3v256x8m81_1 pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D alatch_3v256x8m81_0/ab
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S pmos_1p2$$47337516_3v256x8m81
.ends

.subckt xpredec1_3v256x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1]
+ A[0] clk w_5024_6624# xpredec1_xa_3v256x8m81_7/m3_n46_n5510# vdd vss pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
Xxpredec1_xa_3v256x8m81_0 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[3] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_1 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[1] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_2 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[5] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_3 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[7] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_0 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[0] xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vss vdd xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xxpredec1_xa_3v256x8m81_4 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[2] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_1 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[2] xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vss vdd xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xxpredec1_xa_3v256x8m81_5 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[0] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_2 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[1] xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vss vdd xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_0 vss clk nmos_5p04310591302056_3v256x8m81_1/D vss
+ nmos_5p04310591302056_3v256x8m81
Xxpredec1_xa_3v256x8m81_6 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[4] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_1 nmos_5p04310591302056_3v256x8m81_1/D men vss vss
+ nmos_5p04310591302056_3v256x8m81
Xxpredec1_xa_3v256x8m81_7 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[6] vss xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vdd xpredec1_xa_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 nmos_5p04310591302056_3v256x8m81_1/D xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ vss vss nmos_1p2$$47342636_3v256x8m81
Xpmos_1p2$$47109164_3v256x8m81_0 xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# nmos_5p04310591302056_3v256x8m81_1/D
+ vdd nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81
X0 a_5287_6723# men vdd w_5024_6624# pfet_03v3 ad=0.212p pd=1.46u as=0.5936p ps=3.24u w=1.06u l=0.28u
X1 a_5600_6723# clk nmos_5p04310591302056_3v256x8m81_1/D w_5024_6624# pfet_03v3 ad=0.19345p pd=1.425u as=0.32065p ps=1.665u w=1.06u l=0.28u
X2 nmos_5p04310591302056_3v256x8m81_1/D clk a_5287_6723# w_5024_6624# pfet_03v3 ad=0.32065p pd=1.665u as=0.212p ps=1.46u w=1.06u l=0.28u
X3 vdd men a_5600_6723# w_5024_6624# pfet_03v3 ad=0.5883p pd=3.23u as=0.19345p ps=1.425u w=1.06u l=0.28u
.ends

.subckt pmos_5p04310591302067_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.1196p pd=15.06u as=3.1196p ps=15.06u w=7.09u l=0.28u
.ends

.subckt pmos_1p2$$47643692_3v256x8m81 w_n133_n66# pmos_5p04310591302067_3v256x8m81_0/S
+ pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
Xpmos_5p04310591302067_3v256x8m81_0 pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81
.ends

.subckt nmos_1p2$$47641644_3v256x8m81 nmos_5p04310591302057_3v256x8m81_0/S nmos_5p04310591302057_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v256x8m81_0 nmos_5p04310591302057_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v256x8m81_0/S VSUBS nmos_5p04310591302057_3v256x8m81
.ends

.subckt pmos_1p2$$47642668_3v256x8m81 pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81_0/D
+ a_n14_n34# w_n194_n66#
Xpmos_5p04310591302067_3v256x8m81_0 pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
+ w_n194_n66# pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81
.ends

.subckt xpredec0_xa_3v256x8m81 m3_107_5938# m1_255_3759# a_612_1974# m1_255_3263#
+ m1_255_3619# pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ m1_255_3901# m3_598_2319# pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ a_472_3898# M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
Xpmos_1p2$$47513644_3v256x8m81_0 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_3 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47643692_3v256x8m81_0 pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ a_472_3898# pmos_1p2$$47643692_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_0 nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_1 nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xpmos_1p2$$47642668_3v256x8m81_0 pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S a_612_1974#
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47642668_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_3 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
X0 M3_M2$$47644716_3v256x8m81_2/VSUBS a_612_1974# a_539_2025# M3_M2$$47644716_3v256x8m81_2/VSUBS nfet_03v3 ad=3.1746p pd=12.55u as=1.0439p ps=6.085u w=5.72u l=0.28u
X1 a_539_2025# a_472_3898# pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S M3_M2$$47644716_3v256x8m81_2/VSUBS nfet_03v3 ad=1.0439p pd=6.085u as=3.146p ps=12.54u w=5.72u l=0.28u
.ends

.subckt pmos_5p04310591302063_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.7016p pd=13.16u as=2.7016p ps=13.16u w=6.14u l=0.28u
.ends

.subckt pmos_1p2$$47504428_3v256x8m81 a_n14_n34# pmos_5p04310591302063_3v256x8m81_0/D
+ w_n133_n66# pmos_5p04310591302063_3v256x8m81_0/S
Xpmos_5p04310591302063_3v256x8m81_0 pmos_5p04310591302063_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302063_3v256x8m81_0/S pmos_5p04310591302063_3v256x8m81
.ends

.subckt nmos_5p04310591302065_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.0714p pd=5.75u as=1.0714p ps=5.75u w=2.435u l=0.28u
.ends

.subckt nmos_1p2$$47502380_3v256x8m81 nmos_5p04310591302065_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302065_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302065_3v256x8m81_0 nmos_5p04310591302065_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302065_3v256x8m81_0/S VSUBS nmos_5p04310591302065_3v256x8m81
.ends

.subckt pmos_5p04310591302064_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.6322p pd=17.39u as=3.6322p ps=17.39u w=8.255u l=0.28u
.ends

.subckt pmos_1p2$$47503404_3v256x8m81 pmos_5p04310591302064_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302064_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302064_3v256x8m81_0 pmos_5p04310591302064_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302064_3v256x8m81_0/S pmos_5p04310591302064_3v256x8m81
.ends

.subckt nmos_5p04310591302066_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.4454p pd=7.45u as=1.4454p ps=7.45u w=3.285u l=0.28u
.ends

.subckt xpredec0_bot_3v256x8m81 nmos_5p04310591302066_3v256x8m81_0/D alatch_3v256x8m81_0/a
+ nmos_1p2$$47502380_3v256x8m81_0/nmos_5p04310591302065_3v256x8m81_0/S pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ m1_n74_3354# m1_n74_3071# m1_n74_3213# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/vss
+ m1_n74_2930# m2_800_2096# alatch_3v256x8m81_0/enb pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/S
Xpmos_1p2$$47504428_3v256x8m81_0 nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/S
+ pmos_1p2$$47504428_3v256x8m81
Xnmos_1p2$$47502380_3v256x8m81_0 nmos_1p2$$47502380_3v256x8m81_0/nmos_5p04310591302065_3v256x8m81_0/S
+ nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ alatch_3v256x8m81_0/vss nmos_1p2$$47502380_3v256x8m81
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/enb alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab
+ alatch_3v256x8m81_0/a m2_800_2096# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/vss
+ alatch_3v256x8m81
Xpmos_1p2$$47503404_3v256x8m81_0 pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ alatch_3v256x8m81_0/ab nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ pmos_1p2$$47503404_3v256x8m81
Xnmos_5p04310591302066_3v256x8m81_0 nmos_5p04310591302066_3v256x8m81_0/D alatch_3v256x8m81_0/ab
+ alatch_3v256x8m81_0/vss alatch_3v256x8m81_0/vss nmos_5p04310591302066_3v256x8m81
.ends

.subckt pmos_5p04310591302069_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt xpredec0_3v256x8m81 men x[1] x[2] x[3] A[1] clk xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ x[0] A[0] xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ vdd vss
Xxpredec0_xa_3v256x8m81_3 vss xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D x[3] xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D vss vss xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ vdd xpredec0_xa_3v256x8m81
Xxpredec0_bot_3v256x8m81_0 xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ A[0] vss xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ vdd vss xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ a_4073_6932# pmos_5p04310591302069_3v256x8m81_0/D vdd vdd xpredec0_bot_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 a_4073_6932# pmos_5p04310591302069_3v256x8m81_0/D
+ vss vss nmos_1p2$$46563372_3v256x8m81
Xxpredec0_bot_3v256x8m81_1 xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ A[1] vss xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ vdd vss xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ a_4073_6932# pmos_5p04310591302069_3v256x8m81_0/D vdd vdd xpredec0_bot_3v256x8m81
Xxpredec0_xa_3v256x8m81_0 vss xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D x[0] xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ vss vss xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ vdd xpredec0_xa_3v256x8m81
Xxpredec0_xa_3v256x8m81_1 vss xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D x[2] xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D vss vss xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ vdd xpredec0_xa_3v256x8m81
Xpmos_5p04310591302069_3v256x8m81_0 pmos_5p04310591302069_3v256x8m81_0/D a_4073_6932#
+ a_4073_6932# vdd vdd pmos_5p04310591302069_3v256x8m81
Xxpredec0_xa_3v256x8m81_2 vss xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D x[1] xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ vss vss xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ vdd xpredec0_xa_3v256x8m81
X0 vdd men a_3416_6773# vdd pfet_03v3 ad=0.448p pd=2.72u as=0.162p ps=1.205u w=0.8u l=0.28u
X1 vss clk a_4073_6932# vss nfet_03v3 ad=0.2794p pd=2.15u as=0.1651p ps=1.155u w=0.635u l=0.28u
X2 a_4073_6932# men vss vss nfet_03v3 ad=0.1651p pd=1.155u as=0.2794p ps=2.15u w=0.635u l=0.28u
X3 a_4073_6932# clk a_3091_6773# vdd pfet_03v3 ad=0.218p pd=1.345u as=0.208p ps=1.32u w=0.8u l=0.28u
X4 a_3091_6773# men vdd vdd pfet_03v3 ad=0.208p pd=1.32u as=0.364p ps=2.51u w=0.8u l=0.28u
X5 a_3416_6773# clk a_4073_6932# vdd pfet_03v3 ad=0.162p pd=1.205u as=0.218p ps=1.345u w=0.8u l=0.28u
.ends

.subckt prexdec_top_3v256x8m81 A[2] A[6] xb[3] xc[0] xc[1] xc[2] xb[1] xb[2] xb[0]
+ xa[1] xa[2] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[1] xa[0] xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xa[3] xpredec1_3v256x8m81_0/clk xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/w_5024_6624# xc[3] xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ A[4] men A[5] xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ xpredec0_3v256x8m81_1/clk VSUBS xpredec1_3v256x8m81_0/vdd
Xxpredec1_3v256x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] xpredec1_3v256x8m81_0/clk xpredec1_3v256x8m81_0/w_5024_6624# xpredec1_3v256x8m81_0/vdd
+ xpredec1_3v256x8m81_0/vdd VSUBS xpredec1_3v256x8m81_0/pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd xpredec1_3v256x8m81
Xxpredec0_3v256x8m81_0 men xb[1] xb[2] xb[3] A[4] xpredec0_3v256x8m81_1/clk xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xb[0] A[3] xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/vdd VSUBS xpredec0_3v256x8m81
Xxpredec0_3v256x8m81_1 men xc[1] xc[2] xc[3] A[6] xpredec0_3v256x8m81_1/clk xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xc[0] A[5] xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/vdd VSUBS xpredec0_3v256x8m81
.ends

.subckt pmos_5p04310591302088_3v256x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=2.5608p ps=12.52u w=5.82u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=2.5608p pd=12.52u as=1.5132p ps=6.34u w=5.82u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
.ends

.subckt nmos_5p04310591302081_3v256x8m81 D a_634_n44# a_n168_n44# a_313_n44# a_795_n44#
+ a_474_n44# a_n8_n44# S a_153_n44# VSUBS
X0 D a_153_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X1 D a_474_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X2 D a_n168_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.28u
X3 S a_n8_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X4 D a_795_n44# S VSUBS nfet_03v3 ad=0.1826p pd=1.71u as=0.10892p ps=0.94u w=0.415u l=0.28u
X5 S a_313_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X6 S a_634_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
.ends

.subckt pmos_5p04310591302077_3v256x8m81 D a_n252_n44# a_550_n44# a_229_n44# w_n426_n86#
+ a_390_n44# S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44#
X0 D a_390_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X1 D a_n252_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.968p ps=5.28u w=2.2u l=0.28u
X2 D a_69_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X3 S a_229_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X4 S a_550_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X5 S a_1192_n44# D w_n426_n86# pfet_03v3 ad=0.968p pd=5.28u as=0.572p ps=2.72u w=2.2u l=0.28u
X6 D a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X7 S a_n92_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X9 D a_711_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
.ends

.subckt nmos_5p04310591302075_3v256x8m81 D a_n252_n44# a_550_n44# a_229_n44# a_390_n44#
+ S a_n92_n44# a_1032_n44# a_1192_n44# a_711_n44# a_69_n44# a_871_n44# VSUBS
X0 D a_390_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X1 D a_n252_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.3938p ps=2.67u w=0.895u l=0.28u
X2 D a_69_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X3 S a_229_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X4 S a_550_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X5 S a_1192_n44# D VSUBS nfet_03v3 ad=0.3938p pd=2.67u as=0.2327p ps=1.415u w=0.895u l=0.28u
X6 D a_1032_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X7 S a_n92_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X8 S a_871_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X9 D a_711_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
.ends

.subckt pmos_5p04310591302080_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_5p04310591302076_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt pmos_5p04310591302079_3v256x8m81 D a_486_n44# a_165_n44# a_n156_n44# S a_4_n44#
+ a_646_n44# w_n330_n86# a_808_n44# a_325_n44#
X0 S a_646_n44# D w_n330_n86# pfet_03v3 ad=0.27162p pd=1.555u as=0.2665p ps=1.545u w=1.025u l=0.28u
X1 D a_165_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X2 D a_486_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X3 S a_4_n44# D w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X4 D a_n156_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.451p ps=2.93u w=1.025u l=0.28u
X5 S a_325_n44# D w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X6 D a_808_n44# S w_n330_n86# pfet_03v3 ad=0.451p pd=2.93u as=0.27162p ps=1.555u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302082_3v256x8m81 a_20_n44# D a_181_n44# a_502_n44# a_662_n44#
+ a_n140_n44# S a_341_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X1 S a_662_n44# D w_n314_n86# pfet_03v3 ad=0.5082p pd=3.19u as=0.3003p ps=1.675u w=1.155u l=0.28u
X2 D a_502_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X3 S a_20_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X4 D a_181_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X5 D a_n140_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.5082p ps=3.19u w=1.155u l=0.28u
.ends

.subckt nmos_5p04310591302078_3v256x8m81 D S a_217_n44# a_n104_n44# a_56_n44# VSUBS
X0 D a_217_n44# S VSUBS nfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 S a_56_n44# D VSUBS nfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
X2 D a_n104_n44# S VSUBS nfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
.ends

.subckt wen_v2_3v256x8m81 IGWEN clk wen GWE vss vdd
Xnmos_1p2$$202596396_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_2/S pmos_5p04310591302041_3v256x8m81_1/D
+ vss vss nmos_1p2$$202596396_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_4/D
+ vdd pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_1 pmos_5p04310591302041_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_1/D
+ vdd pmos_5p04310591302041_3v256x8m81_1/S pmos_5p04310591302041_3v256x8m81
Xnmos_5p04310591302081_3v256x8m81_0 pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81_0/S vss pmos_5p04310591302041_3v256x8m81_0/S
+ vss nmos_5p04310591302081_3v256x8m81
Xpmos_5p04310591302077_3v256x8m81_0 IGWEN pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D vdd pmos_5p04310591302082_3v256x8m81_0/D vdd
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302077_3v256x8m81
Xpmos_5p04310591302077_3v256x8m81_2 GWE pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D vdd pmos_5p04310591302079_3v256x8m81_0/D vdd
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302077_3v256x8m81
Xnmos_5p04310591302075_3v256x8m81_0 GWE pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D vss pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D vss nmos_5p04310591302075_3v256x8m81
Xnmos_5p04310591302075_3v256x8m81_1 IGWEN pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D vss pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D vss nmos_5p04310591302075_3v256x8m81
Xpmos_5p04310591302080_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81_2/S vdd vdd pmos_5p04310591302080_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_1/S pmos_5p04310591302014_3v256x8m81_1/D
+ pmos_5p04310591302014_3v256x8m81_3/S vss nmos_5p04310591302010_3v256x8m81
Xnmos_5p04310591302076_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81_2/S vss vss nmos_5p04310591302076_3v256x8m81
Xpmos_1p2$$202587180_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_3/S pmos_5p04310591302014_3v256x8m81_4/D
+ pmos_5p04310591302041_3v256x8m81_1/S vdd pmos_1p2$$202587180_3v256x8m81
Xpmos_5p04310591302079_3v256x8m81_0 pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81_0/S vdd pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S vdd pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_5p04310591302079_3v256x8m81
Xnmos_5p04310591302039_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_4/D
+ pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302041_3v256x8m81_0/S vss nmos_5p04310591302039_3v256x8m81
Xpmos_5p04310591302020_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_1/D
+ pmos_5p04310591302014_3v256x8m81_1/D vdd pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302020_3v256x8m81
Xpmos_1p2$$202586156_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_2/S
+ vdd vdd pmos_1p2$$202586156_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_1/S pmos_5p04310591302014_3v256x8m81_2/S
+ vss vss nmos_1p2$$202595372_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_1 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302041_3v256x8m81_1/S
+ pmos_5p04310591302041_3v256x8m81_1/D vss nmos_1p2$$202595372_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 vdd pmos_5p04310591302079_3v256x8m81_0/D vdd pmos_5p04310591302041_3v256x8m81_0/D
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302082_3v256x8m81_0 wen pmos_5p04310591302082_3v256x8m81_0/D wen wen
+ wen wen vdd wen vdd pmos_5p04310591302082_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_1 pmos_5p04310591302014_3v256x8m81_1/D clk vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_2 vdd pmos_5p04310591302041_3v256x8m81_1/S vdd pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_3 vdd wen vdd pmos_5p04310591302014_3v256x8m81_3/S
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_4 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302014_3v256x8m81_1/D
+ vdd vdd pmos_5p04310591302014_3v256x8m81
Xnmos_5p04310591302078_3v256x8m81_0 pmos_5p04310591302082_3v256x8m81_0/D vss wen wen
+ wen vss nmos_5p04310591302078_3v256x8m81
X0 pmos_5p04310591302014_3v256x8m81_4/D pmos_5p04310591302014_3v256x8m81_1/D vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 vss wen pmos_5p04310591302014_3v256x8m81_3/S vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X2 pmos_5p04310591302014_3v256x8m81_1/D clk vss vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
X3 pmos_5p04310591302041_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_1/D pmos_5p04310591302041_3v256x8m81_0/S vss nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X4 vss pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302041_3v256x8m81_0/D vss nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt nmos_1p2$$48629804_3v256x8m81 nmos_5p04310591302039_3v256x8m81_0/D a_118_n34#
+ a_n41_n34# nmos_5p04310591302039_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302039_3v256x8m81_0 nmos_5p04310591302039_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302039_3v256x8m81_0/S VSUBS nmos_5p04310591302039_3v256x8m81
.ends

.subckt pmos_5p04310591302087_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.6552p pd=22.04u as=4.6552p ps=22.04u w=10.58u l=0.28u
.ends

.subckt pmos_1p2$$47815724_3v256x8m81 pmos_5p04310591302087_3v256x8m81_0/D a_n14_n34#
+ pmos_5p04310591302087_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302087_3v256x8m81_0 pmos_5p04310591302087_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302087_3v256x8m81_0/S pmos_5p04310591302087_3v256x8m81
.ends

.subckt nmos_5p04310591302084_3v256x8m81 a_1394_n44# D a_2357_n44# a_1073_n44# a_2036_n44#
+ a_n51_n44# a_1715_n44# a_752_n44# a_n532_n44# a_431_n44# a_1554_n44# a_591_n44#
+ a_2197_n44# a_n211_n44# S a_110_n44# a_1876_n44# a_1233_n44# a_270_n44# a_912_n44#
+ a_2518_n44# a_n372_n44# VSUBS
X0 S a_270_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X1 D a_1715_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.90167p ps=3.96u w=3.435u l=0.28u
X2 D a_110_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X3 D a_2036_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X4 S a_n51_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X5 S a_591_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X6 D a_1073_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X7 D a_431_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X8 D a_2357_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X9 D a_1394_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X10 S a_n372_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X11 D a_752_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X12 S a_2518_n44# D VSUBS nfet_03v3 ad=1.5114p pd=7.75u as=0.90167p ps=3.96u w=3.435u l=0.28u
X13 S a_1233_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X14 S a_1876_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X15 D a_n211_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X16 S a_2197_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X17 S a_1554_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X18 D a_n532_n44# S VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=1.5114p ps=7.75u w=3.435u l=0.28u
X19 S a_912_n44# D VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
.ends

.subckt nmos_1p2$$48308268_3v256x8m81 nmos_5p04310591302084_3v256x8m81_0/a_752_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1073_n44# nmos_5p04310591302084_3v256x8m81_0/D
+ nmos_5p04310591302084_3v256x8m81_0/a_2036_n44# nmos_5p04310591302084_3v256x8m81_0/a_431_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1715_n44# nmos_5p04310591302084_3v256x8m81_0/a_591_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n532_n44# nmos_5p04310591302084_3v256x8m81_0/a_110_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_270_n44# nmos_5p04310591302084_3v256x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_2197_n44# nmos_5p04310591302084_3v256x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_912_n44# nmos_5p04310591302084_3v256x8m81_0/a_1233_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1876_n44# nmos_5p04310591302084_3v256x8m81_0/S
+ nmos_5p04310591302084_3v256x8m81_0/a_2518_n44# nmos_5p04310591302084_3v256x8m81_0/a_n372_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1394_n44# nmos_5p04310591302084_3v256x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n51_n44# VSUBS
Xnmos_5p04310591302084_3v256x8m81_0 nmos_5p04310591302084_3v256x8m81_0/a_1394_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D nmos_5p04310591302084_3v256x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1073_n44# nmos_5p04310591302084_3v256x8m81_0/a_2036_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n51_n44# nmos_5p04310591302084_3v256x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_752_n44# nmos_5p04310591302084_3v256x8m81_0/a_n532_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_431_n44# nmos_5p04310591302084_3v256x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_591_n44# nmos_5p04310591302084_3v256x8m81_0/a_2197_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n211_n44# nmos_5p04310591302084_3v256x8m81_0/S
+ nmos_5p04310591302084_3v256x8m81_0/a_110_n44# nmos_5p04310591302084_3v256x8m81_0/a_1876_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1233_n44# nmos_5p04310591302084_3v256x8m81_0/a_270_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_912_n44# nmos_5p04310591302084_3v256x8m81_0/a_2518_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n372_n44# VSUBS nmos_5p04310591302084_3v256x8m81
.ends

.subckt nmos_5p04310591302093_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.56u
.ends

.subckt pmos_1p2$$47330348_3v256x8m81 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ pmos_5p04310591302041_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
.ends

.subckt pmos_5p04310591302089_3v256x8m81 a_2502_n44# a_1699_n44# D a_n67_n44# a_2341_n44#
+ a_1378_n44# a_2020_n44# a_1057_n44# a_n548_n44# a_94_n44# a_736_n44# a_n227_n44#
+ a_896_n44# w_n722_n86# S a_415_n44# a_2181_n44# a_1538_n44# a_575_n44# a_1860_n44#
+ a_1217_n44# a_n388_n44# a_254_n44#
X0 D a_n548_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=3.7708p ps=18.02u w=8.57u l=0.28u
X1 S a_575_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X2 D a_415_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X3 D a_1057_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X4 D a_2020_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X5 S a_896_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X6 D a_736_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X7 D a_1378_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X8 D a_2341_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X9 S a_n67_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X10 D a_1699_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.24962p ps=9.095u w=8.57u l=0.28u
X11 S a_2502_n44# D w_n722_n86# pfet_03v3 ad=3.7708p pd=18.02u as=2.24962p ps=9.095u w=8.57u l=0.28u
X12 S a_n388_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X13 S a_1217_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X14 S a_1860_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X15 S a_1538_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X16 S a_2181_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X17 D a_94_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X18 D a_n227_n44# S w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X19 S a_254_n44# D w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
.ends

.subckt pmos_5p04310591302073_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4563p pd=2.275u as=0.7722p ps=4.39u w=1.755u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7722p pd=4.39u as=0.4563p ps=2.275u w=1.755u l=0.28u
.ends

.subckt pmos_1p2$$48623660_3v256x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302073_3v256x8m81_0/D
+ a_118_n34# pmos_5p04310591302073_3v256x8m81_0/S
Xpmos_5p04310591302073_3v256x8m81_0 pmos_5p04310591302073_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302073_3v256x8m81_0/S pmos_5p04310591302073_3v256x8m81
.ends

.subckt pmos_5p04310591302092_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.465u
.ends

.subckt pmos_5p04310591302091_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.004p pd=19.08u as=4.004p ps=19.08u w=9.1u l=0.28u
.ends

.subckt pmos_1p2$$48624684_3v256x8m81 pmos_5p04310591302091_3v256x8m81_0/D a_n14_n34#
+ pmos_5p04310591302091_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302091_3v256x8m81_0 pmos_5p04310591302091_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302091_3v256x8m81_0/S pmos_5p04310591302091_3v256x8m81
.ends

.subckt nmos_5p04310591302083_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1646p pd=1.64u as=0.1646p ps=1.64u w=0.35u l=0.28u
.ends

.subckt nmos_5p04310591302090_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.465u
.ends

.subckt pmos_5p04310591302074_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.56u
.ends

.subckt nmos_5p04310591302085_3v256x8m81 a_530_n44# D a_n112_n44# a_209_n44# a_369_n44#
+ a_48_n44# S VSUBS
X0 D a_n112_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=2.0482p ps=10.19u w=4.655u l=0.28u
X1 S a_369_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=1.22192p ps=5.18u w=4.655u l=0.28u
X3 D a_530_n44# S VSUBS nfet_03v3 ad=2.0482p pd=10.19u as=1.22192p ps=5.18u w=4.655u l=0.28u
X4 S a_48_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
.ends

.subckt nmos_1p2$$48306220_3v256x8m81 a_195_n34# a_n125_n34# a_355_n34# a_34_n34#
+ nmos_5p04310591302085_3v256x8m81_0/D nmos_5p04310591302085_3v256x8m81_0/S VSUBS
+ a_516_n34#
Xnmos_5p04310591302085_3v256x8m81_0 a_516_n34# nmos_5p04310591302085_3v256x8m81_0/D
+ a_n125_n34# a_195_n34# a_355_n34# a_34_n34# nmos_5p04310591302085_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302085_3v256x8m81
.ends

.subckt pmos_5p04310591302094_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3872p pd=2.64u as=0.3872p ps=2.64u w=0.88u l=0.28u
.ends

.subckt nmos_5p04310591302086_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6182p pd=3.69u as=0.6182p ps=3.69u w=1.405u l=0.28u
.ends

.subckt nmos_1p2$$48302124_3v256x8m81 nmos_5p04310591302086_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302086_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302086_3v256x8m81_0 nmos_5p04310591302086_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302086_3v256x8m81_0/S VSUBS nmos_5p04310591302086_3v256x8m81
.ends

.subckt gen_3v256x8_3v256x8m81 VSS tblhl IGWEN cen clk WEN GWE men pmos_5p04310591302088_3v256x8m81_0/D
+ VDD wen_v2_3v256x8m81_0/wen
Xpmos_5p04310591302088_3v256x8m81_0 pmos_5p04310591302088_3v256x8m81_0/D pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ VDD pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_5p04310591302088_3v256x8m81
Xwen_v2_3v256x8m81_0 IGWEN clk wen_v2_3v256x8m81_0/wen GWE VSS VDD wen_v2_3v256x8m81
Xnmos_1p2$$48629804_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S VSS VSS nmos_1p2$$48629804_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_0 VDD tblhl pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ VDD pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_1 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD VDD pmos_1p2$$47815724_3v256x8m81
Xnmos_1p2$$48308268_3v256x8m81_0 pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ men pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D VSS pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ VSS nmos_1p2$$48308268_3v256x8m81
Xnmos_5p04310591302093_3v256x8m81_0 pmos_5p04310591302074_3v256x8m81_0/D clk VSS VSS
+ nmos_5p04310591302093_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_2 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ tblhl VDD VDD pmos_1p2$$47815724_3v256x8m81
Xnmos_5p04310591302093_3v256x8m81_1 pmos_5p04310591302074_3v256x8m81_1/D pmos_5p04310591302074_3v256x8m81_0/D
+ VSS VSS nmos_5p04310591302093_3v256x8m81
Xpmos_1p2$$47330348_3v256x8m81_0 pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ a_3546_5289# pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ VDD pmos_1p2$$47330348_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_3 VDD pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VDD pmos_1p2$$47815724_3v256x8m81
Xpmos_5p04310591302089_3v256x8m81_0 pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ men pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D VDD VDD pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302089_3v256x8m81
Xpmos_1p2$$48623660_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D VDD pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D
+ pmos_5p04310591302094_3v256x8m81_0/D VDD pmos_1p2$$48623660_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_4 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VDD VDD pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_5 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S VDD VDD pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_6 VDD pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_7 VDD pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD pmos_1p2$$47815724_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 clk VSS a_3546_5289# VSS nmos_1p2$$47342636_3v256x8m81
Xpmos_5p04310591302092_3v256x8m81_0 pmos_5p04310591302092_3v256x8m81_0/D pmos_5p04310591302074_3v256x8m81_1/D
+ VDD VDD pmos_5p04310591302092_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_1 men a_3546_5289# VSS VSS nmos_1p2$$47342636_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_0 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_5p04310591302051_3v256x8m81_0/D VDD VDD pmos_1p2$$48624684_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_1 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D VDD VDD pmos_1p2$$48624684_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_0 VDD pmos_5p04310591302051_3v256x8m81_0/D VDD pmos_5p04310591302051_3v256x8m81_0/D
+ pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D pmos_1p2$$46273580_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_2 VDD clk pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ VDD pmos_1p2$$48624684_3v256x8m81
Xnmos_5p04310591302083_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D pmos_5p04310591302092_3v256x8m81_0/D
+ VSS VSS nmos_5p04310591302083_3v256x8m81
Xnmos_5p04310591302090_3v256x8m81_0 pmos_5p04310591302092_3v256x8m81_0/D pmos_5p04310591302074_3v256x8m81_1/D
+ VSS VSS nmos_5p04310591302090_3v256x8m81
Xpmos_5p04310591302074_3v256x8m81_0 pmos_5p04310591302074_3v256x8m81_0/D clk VDD VDD
+ pmos_5p04310591302074_3v256x8m81
Xpmos_5p04310591302074_3v256x8m81_1 pmos_5p04310591302074_3v256x8m81_1/D pmos_5p04310591302074_3v256x8m81_0/D
+ VDD VDD pmos_5p04310591302074_3v256x8m81
Xnmos_1p2$$48306220_3v256x8m81_0 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_5p04310591302088_3v256x8m81_0/D
+ VSS VSS pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S nmos_1p2$$48306220_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S VDD VDD pmos_5p04310591302051_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 a_3546_5289# VSS pmos_1p2$$46285868_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_5p04310591302094_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D pmos_5p04310591302092_3v256x8m81_0/D
+ VDD VDD pmos_5p04310591302094_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_1 pmos_5p04310591302051_3v256x8m81_0/D pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ VSS VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 VDD VDD pmos_1p2$$46285868_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ a_3546_5289# pmos_1p2$$46285868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 cen a_3546_5289# pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ VSS nmos_1p2$$46551084_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_2 pmos_1p2$$46285868_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D
+ pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_1 VDD pmos_1p2$$47330348_3v256x8m81_0/pmos_5p04310591302041_3v256x8m81_0/S
+ cen pmos_1p2$$46285868_3v256x8m81_0/pmos_5p04310591302014_3v256x8m81_0/D pmos_1p2$$46285868_3v256x8m81
Xnmos_1p2$$48302124_3v256x8m81_0 VSS pmos_5p04310591302094_3v256x8m81_0/D pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D
+ VSS nmos_1p2$$48302124_3v256x8m81
X0 a_8790_2243# tblhl pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X1 a_3606_4291# men VDD VDD pfet_03v3 ad=0.2769p pd=1.585u as=0.50587p ps=3.08u w=1.065u l=0.28u
X2 a_7891_338# pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X3 a_6888_183# clk a_6728_183# VSS nfet_03v3 ad=2.7521p pd=11.105u as=2.7521p ps=11.105u w=10.585u l=0.28u
X4 VSS pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S a_7891_338# VSS nfet_03v3 ad=3.93622p pd=17.86u as=2.2009p ps=8.985u w=8.465u l=0.28u
X5 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S tblhl a_8470_2243# VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X6 a_8470_2243# pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VSS VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.96232p ps=5.14u w=2.115u l=0.28u
X7 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S pmos_5p04310591302051_3v256x8m81_0/D a_6888_183# VSS nfet_03v3 ad=5.2925p pd=22.17u as=2.7521p ps=11.105u w=10.585u l=0.28u
X8 a_7571_338# pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VSS VSS nfet_03v3 ad=2.2009p pd=8.985u as=3.85157p ps=17.84u w=8.465u l=0.28u
X9 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S a_7571_338# VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X10 a_6728_183# pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D VSS VSS nfet_03v3 ad=2.7521p pd=11.105u as=4.6574p ps=22.05u w=10.585u l=0.28u
X11 a_3546_5289# clk a_3606_4291# VDD pfet_03v3 ad=0.50587p pd=3.08u as=0.2769p ps=1.585u w=1.065u l=0.28u
X12 VSS pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S a_8790_2243# VSS nfet_03v3 ad=0.99405p pd=5.17u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt control_3v256x8_3v256x8m81 RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[2] A[0] xb[1] xc[3] xc[1] xc[2] xa[1] A[9]
+ A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWE GWEN ypredec1_3v256x8m81_0/ly[1]
+ ypredec1_3v256x8m81_0/ly[2] ypredec1_3v256x8m81_0/ly[4] xa[3] ypredec1_3v256x8m81_0/ly[5]
+ ypredec1_3v256x8m81_0/ly[6] xa[0] ypredec1_3v256x8m81_0/ly[7] CEN xc[0] men prexdec_top_3v256x8m81_0/xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ VSS VDD
Xypredec1_3v256x8m81_0 ypredec1_3v256x8m81_0/ly[5] ypredec1_3v256x8m81_0/ly[4] ypredec1_3v256x8m81_0/ly[7]
+ ypredec1_3v256x8m81_0/ly[2] ypredec1_3v256x8m81_0/ly[1] LYS[7] RYS[0] RYS[1] RYS[2]
+ RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_3v256x8m81_0/ly[6] men A[0] A[1] A[2]
+ CLK A[1] VDD A[0] VDD A[2] VDD VDD VDD VSS VDD ypredec1_3v256x8m81
Xprexdec_top_3v256x8m81_0 A[5] A[9] xb[3] xc[0] xc[1] xc[2] xb[1] xb[2] xb[0] xa[1]
+ xa[2] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[4] xa[0] VSS xa[3] CLK VSS VSS VDD xc[3]
+ VSS VDD A[7] men A[8] prexdec_top_3v256x8m81_0/xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ CLK VSS VDD prexdec_top_3v256x8m81
Xgen_3v256x8_3v256x8m81_0 VSS tblhl IGWEN CEN CLK gen_3v256x8_3v256x8m81_0/WEN GWE
+ men gen_3v256x8_3v256x8m81_0/pmos_5p04310591302088_3v256x8m81_0/D VDD GWEN gen_3v256x8_3v256x8m81
.ends

.subckt pmos_5p043105913020101_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_5p043105913020107_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.6058p pd=2.85u as=1.0252p ps=5.54u w=2.33u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=1.0252p pd=5.54u as=0.6058p ps=2.85u w=2.33u l=0.28u
.ends

.subckt pmos_5p043105913020103_3v256x8m81 D a_265_n44# S a_n56_n44# a_104_n44# w_n230_n86#
X0 D a_265_n44# S w_n230_n86# pfet_03v3 ad=2.0526p pd=10.21u as=1.22455p ps=5.19u w=4.665u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=1.2129p pd=5.185u as=2.0526p ps=10.21u w=4.665u l=0.28u
X2 S a_104_n44# D w_n230_n86# pfet_03v3 ad=1.22455p pd=5.19u as=1.2129p ps=5.185u w=4.665u l=0.28u
.ends

.subckt pmos_1p2_03_R270_3v256x8m81 a_n69_n138# pmos_5p043105913020103_3v256x8m81_0/S
+ a_90_n138# w_n138_n63# a_251_n138# pmos_5p043105913020103_3v256x8m81_0/D
Xpmos_5p043105913020103_3v256x8m81_0 pmos_5p043105913020103_3v256x8m81_0/D a_251_n138#
+ pmos_5p043105913020103_3v256x8m81_0/S a_n69_n138# a_90_n138# w_n138_n63# pmos_5p043105913020103_3v256x8m81
.ends

.subckt pmos_5p043105913020108_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6669p pd=3.085u as=1.1286p ps=6.01u w=2.565u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1286p pd=6.01u as=0.6669p ps=3.085u w=2.565u l=0.28u
.ends

.subckt pmos_1p2_01_R270_3v256x8m81 pmos_5p043105913020108_3v256x8m81_0/D w_n246_n93#
+ a_118_n33# pmos_5p043105913020108_3v256x8m81_0/S a_n41_n33#
Xpmos_5p043105913020108_3v256x8m81_0 pmos_5p043105913020108_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n246_n93# pmos_5p043105913020108_3v256x8m81_0/S pmos_5p043105913020108_3v256x8m81
.ends

.subckt nmos_1p2_02_R270_3v256x8m81 nmos_5p04310591302044_3v256x8m81_0/S a_n14_n33#
+ nmos_5p04310591302044_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302044_3v256x8m81_0 nmos_5p04310591302044_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302044_3v256x8m81_0/S VSUBS nmos_5p04310591302044_3v256x8m81
.ends

.subckt nmos_5p043105913020109_3v256x8m81 D a_n28_n44# a_132_n44# S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S a_132_n44# D VSUBS nfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_5p043105913020110_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3256p pd=2.36u as=0.3256p ps=2.36u w=0.74u l=0.28u
.ends

.subckt pmos_5p043105913020104_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_1p2_02_R270_3v256x8m81 a_118_n33# a_n41_n33# pmos_5p043105913020104_3v256x8m81_0/D
+ w_n138_n63# pmos_5p043105913020104_3v256x8m81_0/S
Xpmos_5p043105913020104_3v256x8m81_0 pmos_5p043105913020104_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020104_3v256x8m81_0/S pmos_5p043105913020104_3v256x8m81
.ends

.subckt nmos_5p043105913020106_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1601p pd=1.64u as=0.1601p ps=1.64u w=0.305u l=0.28u
.ends

.subckt pmos_5p043105913020105_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.28u
.ends

.subckt xdec_3v256x8m81 RWL LWL men xc xb xa m2_11898_n156# m2_9070_n156# m2_7748_n156#
+ m2_8806_n156# m2_10577_n156# m2_10840_n156# m2_7219_n156# m2_7483_n156# m2_11634_n156#
+ m2_12427_n156# m2_8277_n156# m2_8541_n156# m2_11105_n156# vss m2_11370_n156# m2_12163_n156#
+ m2_8012_n156# vdd
Xnmos_5p043105913020107_3v256x8m81_0 LWL pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vss vss nmos_5p043105913020107_3v256x8m81
Xpmos_1p2_03_R270_3v256x8m81_0 pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ LWL pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vdd pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd pmos_1p2_03_R270_3v256x8m81
Xnmos_5p043105913020107_3v256x8m81_1 RWL pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D vss vss nmos_5p043105913020107_3v256x8m81
Xpmos_1p2_01_R270_3v256x8m81_0 pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd nmos_5p043105913020109_3v256x8m81_0/S vdd nmos_5p043105913020109_3v256x8m81_0/S
+ pmos_1p2_01_R270_3v256x8m81
Xpmos_1p2_01_R270_3v256x8m81_1 pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd nmos_5p043105913020109_3v256x8m81_0/S vdd nmos_5p043105913020109_3v256x8m81_0/S
+ pmos_1p2_01_R270_3v256x8m81
Xnmos_1p2_02_R270_3v256x8m81_0 nmos_5p043105913020109_3v256x8m81_0/S pmos_5p043105913020105_3v256x8m81_3/S
+ vss vss nmos_1p2_02_R270_3v256x8m81
Xnmos_5p043105913020109_3v256x8m81_0 men pmos_5p043105913020110_3v256x8m81_0/S pmos_5p043105913020110_3v256x8m81_0/S
+ nmos_5p043105913020109_3v256x8m81_0/S vss nmos_5p043105913020109_3v256x8m81
Xpmos_5p043105913020103_3v256x8m81_0 vdd pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ RWL pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd pmos_5p043105913020103_3v256x8m81
Xpmos_5p043105913020110_3v256x8m81_0 vdd pmos_5p043105913020105_3v256x8m81_3/S vdd
+ pmos_5p043105913020110_3v256x8m81_0/S pmos_5p043105913020110_3v256x8m81
Xpmos_1p2_02_R270_3v256x8m81_0 pmos_5p043105913020105_3v256x8m81_3/S pmos_5p043105913020105_3v256x8m81_3/S
+ men vdd nmos_5p043105913020109_3v256x8m81_0/S pmos_1p2_02_R270_3v256x8m81
Xnmos_5p043105913020106_3v256x8m81_0 vss pmos_5p043105913020105_3v256x8m81_3/S pmos_5p043105913020110_3v256x8m81_0/S
+ vss nmos_5p043105913020106_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_1 pmos_5p043105913020105_3v256x8m81_3/S xb vdd
+ vdd pmos_5p043105913020105_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_2 vdd xa vdd pmos_5p043105913020105_3v256x8m81_3/S
+ pmos_5p043105913020105_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_3 vdd xc vdd pmos_5p043105913020105_3v256x8m81_3/S
+ pmos_5p043105913020105_3v256x8m81
X0 vss xc a_9450_422# vss nfet_03v3 ad=0.88935p pd=4.15u as=0.29032p ps=1.865u w=1.47u l=0.28u
X1 vss nmos_5p043105913020109_3v256x8m81_0/S pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vss nfet_03v3 ad=0.2796p pd=4.9u as=1.0252p ps=5.54u w=2.33u l=0.28u
X2 a_9450_280# xa pmos_5p043105913020105_3v256x8m81_3/S vss nfet_03v3 ad=0.31605p pd=1.9u as=0.74235p ps=3.95u w=1.47u l=0.28u
X3 a_9450_422# xb a_9450_280# vss nfet_03v3 ad=0.29032p pd=1.865u as=0.31605p ps=1.9u w=1.47u l=0.28u
X4 vss nmos_5p043105913020109_3v256x8m81_0/S pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D vss nfet_03v3 ad=1.15335p pd=5.65u as=1.0718p ps=5.58u w=2.33u l=0.28u
.ends

.subckt xdec8_3v256x8m81 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] RWL[7] LWL[1] LWL[7]
+ LWL[6] LWL[0] LWL[3] xa[4] xa[7] xa[1] xa[3] xa[0] xa[6] xdec_3v256x8m81_7/m2_10577_n156#
+ RWL[3] xdec_3v256x8m81_7/m2_7219_n156# xb xdec_3v256x8m81_7/m2_11634_n156# xa[5]
+ xa[2] RWL[0] xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_12427_n156# RWL[6]
+ xdec_3v256x8m81_7/m2_11898_n156# xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_10840_n156#
+ men xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8541_n156#
+ xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8277_n156# RWL[1] xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_8012_n156# vss vdd xdec_3v256x8m81_7/m2_11105_n156# xc
Xxdec_3v256x8m81_6 RWL[3] LWL[3] men xc xb xa[3] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_7 RWL[1] LWL[1] men xc xb xa[1] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_0 RWL[6] LWL[6] men xc xb xa[6] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_1 RWL[4] LWL[4] men xc xb xa[4] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_2 RWL[2] LWL[2] men xc xb xa[2] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_3 RWL[0] LWL[0] men xc xb xa[0] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_4 RWL[7] LWL[7] men xc xb xa[7] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
Xxdec_3v256x8m81_5 RWL[5] LWL[5] men xc xb xa[5] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ xdec_3v256x8m81_7/m2_8277_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ vss xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8012_n156#
+ vdd xdec_3v256x8m81
.ends

.subckt xdec32_3v256x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[14] RWL[13] LWL[9] LWL[8]
+ LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[8] RWL[5] RWL[3] RWL[0]
+ RWL[2] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6]
+ LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19]
+ RWL[23] RWL[24] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[7]
+ xb[3] xb[2] xb[0] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156# RWL[20] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[6] RWL[21] RWL[25] xa[3] xa[0] RWL[28] RWL[1] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ RWL[7] xc RWL[4] RWL[16] xa[5] RWL[9] RWL[29] RWL[22] xa[4] xb[1] RWL[15] RWL[26]
+ xa[1] RWL[12] vdd vss
Xxdec8_3v256x8m81_0 LWL[29] LWL[28] LWL[26] RWL[29] RWL[28] RWL[26] RWL[31] LWL[25]
+ LWL[31] LWL[30] LWL[24] LWL[27] xa[4] xa[7] xa[1] xa[3] xa[0] xa[6] xa[7] RWL[27]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156# xb[3] xa[3] xa[5] xa[2] RWL[24]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156# xa[0] RWL[30] xa[2] xb[0] xa[6]
+ men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156# xa[4] xb[2] xa[1] xb[3] RWL[25]
+ xb[1] xc vss vdd xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_1 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] RWL[7] LWL[1] LWL[7]
+ LWL[6] LWL[0] LWL[3] xa[4] xa[7] xa[1] xa[3] xa[0] xa[6] xa[7] RWL[3] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156#
+ xb[0] xa[3] xa[5] xa[2] RWL[0] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[0] RWL[6] xa[2] xb[0] xa[6] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ xa[4] xb[2] xa[1] xb[3] RWL[1] xb[1] xc vss vdd xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_2 LWL[13] LWL[12] LWL[10] RWL[13] RWL[12] RWL[10] RWL[15] LWL[9]
+ LWL[15] LWL[14] LWL[8] LWL[11] xa[4] xa[7] xa[1] xa[3] xa[0] xa[6] xa[7] RWL[11]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156# xb[1] xa[3] xa[5] xa[2] RWL[8]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156# xa[0] RWL[14] xa[2] xb[0] xa[6]
+ men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156# xa[4] xb[2] xa[1] xb[3] RWL[9]
+ xb[1] xc vss vdd xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_3 LWL[21] LWL[20] LWL[18] RWL[21] RWL[20] RWL[18] RWL[23] LWL[17]
+ LWL[23] LWL[22] LWL[16] LWL[19] xa[4] xa[7] xa[1] xa[3] xa[0] xa[6] xa[7] RWL[19]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156# xb[2] xa[3] xa[5] xa[2] RWL[16]
+ xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156# xa[0] RWL[22] xa[2] xb[0] xa[6]
+ men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156# xa[4] xb[2] xa[1] xb[3] RWL[17]
+ xb[1] xc vss vdd xa[5] xc xdec8_3v256x8m81
.ends

.subckt pmos_5p043105913020100_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.5314p pd=6.41u as=2.5916p ps=12.66u w=5.89u l=0.28u
X1 S a_132_n44# D w_n202_n86# pfet_03v3 ad=2.5916p pd=12.66u as=1.5314p ps=6.41u w=5.89u l=0.28u
.ends

.subckt pmos_1p2_02_R90_3v256x8m81 pmos_5p043105913020100_3v256x8m81_0/D w_n138_n63#
+ a_118_n33# pmos_5p043105913020100_3v256x8m81_0/S a_n41_n33#
Xpmos_5p043105913020100_3v256x8m81_0 pmos_5p043105913020100_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020100_3v256x8m81_0/S pmos_5p043105913020100_3v256x8m81
.ends

.subckt nmos_5p04310591302099_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.0746p pd=10.31u as=2.0746p ps=10.31u w=4.715u l=0.28u
.ends

.subckt nmos_5p043105913020111_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.5412p pd=3.34u as=0.5412p ps=3.34u w=1.23u l=0.28u
.ends

.subckt pmoscap_R270_3v256x8m81 m3_770_16# a_n126_928# a_n140_236# m3_152_0# w_n226_n219#
X0 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=1.20555p pd=6.07u as=0 ps=0 w=2.565u l=2.505u
X1 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=0.6733p pd=3.09u as=0 ps=0 w=2.565u l=2.505u
.ends

.subckt nmos_1p2_02_R90_3v256x8m81 nmos_5p04310591302099_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302099_3v256x8m81_0 nmos_5p04310591302099_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v256x8m81_0/S VSUBS nmos_5p04310591302099_3v256x8m81
.ends

.subckt pmoscap_L1_W2_R270_3v256x8m81 m3_307_0# m3_600_0# a_597_236# m1_38_36# M1_NACTIVE_01_R270_3v256x8m81_0/VSUBS
+ a_8_236#
X0 a_597_236# M1_NACTIVE_01_R270_3v256x8m81_0/VSUBS a_8_236# m1_38_36# pfet_03v3 ad=1.1286p pd=6.01u as=1.1286p ps=6.01u w=2.565u l=2.505u
.ends

.subckt nmos_5p043105913020102_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_1p2_01_R270_3v256x8m81 nmos_5p043105913020102_3v256x8m81_0/D a_n14_n33#
+ VSUBS nmos_5p043105913020102_3v256x8m81_0/S
Xnmos_5p043105913020102_3v256x8m81_0 nmos_5p043105913020102_3v256x8m81_0/D a_n14_n33#
+ nmos_5p043105913020102_3v256x8m81_0/S VSUBS nmos_5p043105913020102_3v256x8m81
.ends

.subckt pmos_1p2_01_R90_3v256x8m81 pmos_5p043105913020101_3v256x8m81_0/S w_n137_n63#
+ pmos_5p043105913020101_3v256x8m81_0/D a_n14_n33#
Xpmos_5p043105913020101_3v256x8m81_0 pmos_5p043105913020101_3v256x8m81_0/D a_n14_n33#
+ w_n137_n63# pmos_5p043105913020101_3v256x8m81_0/S pmos_5p043105913020101_3v256x8m81
.ends

.subckt xdec64_3v256x8m81 DRWL DLWL LWL[20] LWL[21] LWL[22] LWL[27] LWL[13] LWL[14]
+ LWL[16] LWL[3] LWL[2] LWL[1] LWL[0] LWL[8] LWL[9] LWL[7] LWL[30] RWL[31] RWL[30]
+ RWL[29] RWL[22] RWL[4] RWL[2] RWL[0] RWL[1] RWL[3] RWL[7] RWL[9] RWL[11] RWL[14]
+ RWL[15] RWL[16] RWL[17] RWL[18] RWL[19] RWL[20] xb[0] xb[1] xb[2] xb[3] xa[7] xa[6]
+ xa[5] xa[4] xa[0] men xa[3] xa[2] xa[1] xc[1] RWL[21] LWL[25] LWL[28] LWL[26] LWL[11]
+ LWL[12] LWL[24] RWL[27] LWL[23] LWL[10] LWL[31] LWL[19] RWL[12] LWL[17] RWL[28]
+ RWL[25] xc[0] RWL[10] LWL[29] RWL[5] RWL[26] vss LWL[5] LWL[6] RWL[13] LWL[18] RWL[24]
+ RWL[8] LWL[4] LWL[15] vdd RWL[23] RWL[6]
Xpmos_5p043105913020101_3v256x8m81_0 vdd pmos_5p043105913020101_3v256x8m81_1/D vdd
+ pmos_5p043105913020101_3v256x8m81_0/S pmos_5p043105913020101_3v256x8m81
Xpmos_5p043105913020101_3v256x8m81_1 pmos_5p043105913020101_3v256x8m81_1/D vss vdd
+ men pmos_5p043105913020101_3v256x8m81
Xxdec32_3v256x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[14] RWL[13] LWL[9] LWL[8] LWL[0]
+ LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[8] RWL[5] RWL[3] RWL[0] RWL[2]
+ LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6] LWL[28]
+ LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19] RWL[23]
+ RWL[24] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[7] xb[3]
+ xb[2] xb[0] vdd RWL[20] vdd xa[6] RWL[21] RWL[25] xa[3] xa[0] RWL[28] RWL[1] men
+ xc[1] RWL[7] xc[0] RWL[4] RWL[16] xa[5] RWL[9] RWL[29] RWL[22] xa[4] xb[1] RWL[15]
+ RWL[26] xa[1] RWL[12] vdd vss xdec32_3v256x8m81
Xpmos_1p2_02_R90_3v256x8m81_0 DLWL vdd nmos_5p043105913020111_3v256x8m81_0/S vdd nmos_5p043105913020111_3v256x8m81_0/S
+ pmos_1p2_02_R90_3v256x8m81
Xpmos_1p2_02_R90_3v256x8m81_1 DRWL vdd pmos_5p043105913020101_3v256x8m81_0/S vdd pmos_5p043105913020101_3v256x8m81_0/S
+ pmos_1p2_02_R90_3v256x8m81
Xnmos_5p04310591302099_3v256x8m81_0 vss pmos_5p043105913020101_3v256x8m81_0/S DRWL
+ vss nmos_5p04310591302099_3v256x8m81
Xnmos_5p043105913020111_3v256x8m81_0 vss pmos_5p043105913020101_3v256x8m81_1/D nmos_5p043105913020111_3v256x8m81_0/S
+ vss nmos_5p043105913020111_3v256x8m81
Xnmos_5p043105913020111_3v256x8m81_1 vss pmos_5p043105913020101_3v256x8m81_1/D pmos_5p043105913020101_3v256x8m81_0/S
+ vss nmos_5p043105913020111_3v256x8m81
Xpmoscap_R270_3v256x8m81_0 RWL[16] vss vdd RWL[17] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_1 RWL[14] vss vdd RWL[15] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_2 RWL[12] vss vdd RWL[13] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_3 RWL[10] vss vdd RWL[11] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_4 RWL[8] vss vdd RWL[9] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_5 RWL[6] vss vdd RWL[7] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_6 RWL[4] vss vdd RWL[5] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_7 RWL[2] vss vdd RWL[3] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_8 RWL[0] vss vdd RWL[1] vdd pmoscap_R270_3v256x8m81
Xnmos_1p2_02_R90_3v256x8m81_0 vss nmos_5p043105913020111_3v256x8m81_0/S DLWL vss nmos_1p2_02_R90_3v256x8m81
Xpmoscap_R270_3v256x8m81_9 RWL[30] vss vdd RWL[31] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_30 LWL[20] vss vdd LWL[21] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_31 LWL[18] vss vdd LWL[19] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_20 LWL[8] vss vdd LWL[9] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_10 RWL[28] vss vdd RWL[29] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_21 LWL[6] vss vdd LWL[7] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_11 RWL[26] vss vdd RWL[27] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_22 LWL[4] vss vdd LWL[5] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_12 RWL[24] vss vdd RWL[25] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_23 LWL[2] vss vdd LWL[3] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_13 RWL[22] vss vdd RWL[23] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_24 LWL[0] vss vdd LWL[1] vdd pmoscap_R270_3v256x8m81
Xpmoscap_L1_W2_R270_3v256x8m81_0 DLWL vdd vdd vdd vss vdd pmoscap_L1_W2_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_25 LWL[30] vss vdd LWL[31] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_14 RWL[20] vss vdd RWL[21] vdd pmoscap_R270_3v256x8m81
Xpmoscap_L1_W2_R270_3v256x8m81_1 DRWL vdd vdd vdd vss vdd pmoscap_L1_W2_R270_3v256x8m81
Xnmos_1p2_01_R270_3v256x8m81_0 men vdd vss pmos_5p043105913020101_3v256x8m81_1/D nmos_1p2_01_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_26 LWL[28] vss vdd LWL[29] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_15 RWL[18] vss vdd RWL[19] vdd pmoscap_R270_3v256x8m81
Xpmos_1p2_01_R90_3v256x8m81_0 nmos_5p043105913020111_3v256x8m81_0/S vdd vdd pmos_5p043105913020101_3v256x8m81_1/D
+ pmos_1p2_01_R90_3v256x8m81
Xpmoscap_R270_3v256x8m81_27 LWL[26] vss vdd LWL[27] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_16 LWL[16] vss vdd LWL[17] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_28 LWL[24] vss vdd LWL[25] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_29 LWL[22] vss vdd LWL[23] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_17 LWL[14] vss vdd LWL[15] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_18 LWL[12] vss vdd LWL[13] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_19 LWL[10] vss vdd LWL[11] vdd pmoscap_R270_3v256x8m81
.ends

.subckt gf180mcu_ocd_ip_sram__sram256x8m8wm1 A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+ CEN CLK D[7] D[5] D[3] D[1] GWEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] VDD WEN[7]
+ WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1] WEN[0] VSS
Xlcol4_256_3v256x8m81_0 lcol4_256_3v256x8m81_0/WL[20] xdec64_3v256x8m81_0/LWL[20]
+ lcol4_256_3v256x8m81_0/WL[18] VSS VSS lcol4_256_3v256x8m81_0/WL[13] VSS VSS xdec64_3v256x8m81_0/LWL[9]
+ lcol4_256_3v256x8m81_0/WL[8] xdec64_3v256x8m81_0/LWL[7] lcol4_256_3v256x8m81_0/WL[6]
+ xdec64_3v256x8m81_0/LWL[5] xdec64_3v256x8m81_0/LWL[4] xdec64_3v256x8m81_0/LWL[3]
+ xdec64_3v256x8m81_0/LWL[2] xdec64_3v256x8m81_0/LWL[1] lcol4_256_3v256x8m81_0/WL[31]
+ lcol4_256_3v256x8m81_0/din[1] lcol4_256_3v256x8m81_0/din[3] lcol4_256_3v256x8m81_0/din[2]
+ lcol4_256_3v256x8m81_0/q[1] lcol4_256_3v256x8m81_0/q[2] lcol4_256_3v256x8m81_0/q[3]
+ lcol4_256_3v256x8m81_0/pcb[2] lcol4_256_3v256x8m81_0/pcb[3] lcol4_256_3v256x8m81_0/pcb[0]
+ lcol4_256_3v256x8m81_0/pcb[1] WEN[0] WEN[1] WEN[2] WEN[3] rcol4_256_3v256x8m81_0/GWE
+ Q[0] Q[1] control_3v256x8_3v256x8m81_0/IGWEN xdec64_3v256x8m81_0/LWL[6] rcol4_256_3v256x8m81_0/GWE
+ xdec64_3v256x8m81_0/LWL[8] xdec64_3v256x8m81_0/LWL[21] D[1] xdec64_3v256x8m81_0/LWL[22]
+ xdec64_3v256x8m81_0/LWL[23] xdec64_3v256x8m81_0/LWL[24] xdec64_3v256x8m81_0/LWL[25]
+ xdec64_3v256x8m81_0/LWL[26] xdec64_3v256x8m81_0/LWL[27] D[3] xdec64_3v256x8m81_0/LWL[28]
+ xdec64_3v256x8m81_0/LWL[29] Q[3] Q[2] control_3v256x8_3v256x8m81_0/LYS[7] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[1]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[2] VDD rcol4_256_3v256x8m81_0/GWE
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[4] xdec64_3v256x8m81_0/men xdec64_3v256x8m81_0/LWL[10]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[5] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[6]
+ xdec64_3v256x8m81_0/LWL[11] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[7]
+ xdec64_3v256x8m81_0/LWL[12] rcol4_256_3v256x8m81_0/GWE xdec64_3v256x8m81_0/LWL[30]
+ xdec64_3v256x8m81_0/LWL[13] xdec64_3v256x8m81_0/LWL[14] xdec64_3v256x8m81_0/LWL[31]
+ xdec64_3v256x8m81_0/LWL[15] xdec64_3v256x8m81_0/LWL[16] xdec64_3v256x8m81_0/LWL[17]
+ xdec64_3v256x8m81_0/LWL[18] rcol4_256_3v256x8m81_0/GWE xdec64_3v256x8m81_0/LWL[0]
+ xdec64_3v256x8m81_0/LWL[19] VSS VDD lcol4_256_3v256x8m81
Xrcol4_256_3v256x8m81_0 xdec64_3v256x8m81_0/RWL[30] rcol4_256_3v256x8m81_0/WL[20]
+ xdec64_3v256x8m81_0/RWL[28] xdec64_3v256x8m81_0/RWL[31] VSS xdec64_3v256x8m81_0/RWL[16]
+ rcol4_256_3v256x8m81_0/WL[31] VSS VSS xdec64_3v256x8m81_0/RWL[27] xdec64_3v256x8m81_0/RWL[20]
+ xdec64_3v256x8m81_0/RWL[29] VSS rcol4_256_3v256x8m81_0/WL[8] xdec64_3v256x8m81_0/RWL[5]
+ VSS rcol4_256_3v256x8m81_0/WL[13] rcol4_256_3v256x8m81_0/WL[6] rcol4_256_3v256x8m81_0/tblhl
+ rcol4_256_3v256x8m81_0/GWE xdec64_3v256x8m81_0/RWL[11] rcol4_256_3v256x8m81_0/din[7]
+ rcol4_256_3v256x8m81_0/q[5] rcol4_256_3v256x8m81_0/q[6] rcol4_256_3v256x8m81_0/q[7]
+ rcol4_256_3v256x8m81_0/din[5] rcol4_256_3v256x8m81_0/din[6] rcol4_256_3v256x8m81_0/q[4]
+ rcol4_256_3v256x8m81_0/pcb[7] rcol4_256_3v256x8m81_0/pcb[4] WEN[7] WEN[4] rcol4_256_3v256x8m81_0/pcb[5]
+ WEN[6] WEN[5] xdec64_3v256x8m81_0/RWL[17] rcol4_256_3v256x8m81_0/saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb
+ xdec64_3v256x8m81_0/RWL[14] xdec64_3v256x8m81_0/RWL[13] control_3v256x8_3v256x8m81_0/RYS[1]
+ xdec64_3v256x8m81_0/men D[7] Q[6] xdec64_3v256x8m81_0/RWL[21] control_3v256x8_3v256x8m81_0/RYS[6]
+ xdec64_3v256x8m81_0/RWL[19] xdec64_3v256x8m81_0/RWL[15] control_3v256x8_3v256x8m81_0/RYS[7]
+ rcol4_256_3v256x8m81_0/saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb control_3v256x8_3v256x8m81_0/RYS[2]
+ xdec64_3v256x8m81_0/RWL[8] xdec64_3v256x8m81_0/RWL[22] xdec64_3v256x8m81_0/RWL[7]
+ xdec64_3v256x8m81_0/RWL[6] xdec64_3v256x8m81_0/RWL[1] xdec64_3v256x8m81_0/RWL[0]
+ control_3v256x8_3v256x8m81_0/RYS[0] xdec64_3v256x8m81_0/DRWL xdec64_3v256x8m81_0/RWL[10]
+ xdec64_3v256x8m81_0/RWL[9] xdec64_3v256x8m81_0/RWL[24] xdec64_3v256x8m81_0/RWL[23]
+ control_3v256x8_3v256x8m81_0/RYS[5] Q[7] Q[4] xdec64_3v256x8m81_0/RWL[2] control_3v256x8_3v256x8m81_0/RYS[4]
+ VSS Q[5] D[5] xdec64_3v256x8m81_0/RWL[12] xdec64_3v256x8m81_0/RWL[26] control_3v256x8_3v256x8m81_0/IGWEN
+ control_3v256x8_3v256x8m81_0/RYS[3] xdec64_3v256x8m81_0/RWL[25] xdec64_3v256x8m81_0/RWL[4]
+ xdec64_3v256x8m81_0/RWL[3] xdec64_3v256x8m81_0/RWL[18] VDD VSS rcol4_256_3v256x8m81
Xcontrol_3v256x8_3v256x8m81_0 control_3v256x8_3v256x8m81_0/RYS[7] control_3v256x8_3v256x8m81_0/RYS[6]
+ control_3v256x8_3v256x8m81_0/RYS[5] control_3v256x8_3v256x8m81_0/RYS[4] control_3v256x8_3v256x8m81_0/RYS[3]
+ control_3v256x8_3v256x8m81_0/RYS[2] control_3v256x8_3v256x8m81_0/RYS[1] control_3v256x8_3v256x8m81_0/RYS[0]
+ VSS control_3v256x8_3v256x8m81_0/LYS[1] control_3v256x8_3v256x8m81_0/LYS[2] control_3v256x8_3v256x8m81_0/LYS[3]
+ control_3v256x8_3v256x8m81_0/LYS[6] control_3v256x8_3v256x8m81_0/LYS[5] control_3v256x8_3v256x8m81_0/LYS[4]
+ control_3v256x8_3v256x8m81_0/LYS[7] rcol4_256_3v256x8m81_0/tblhl control_3v256x8_3v256x8m81_0/IGWEN
+ xdec64_3v256x8m81_0/xb[3] xdec64_3v256x8m81_0/xb[2] xdec64_3v256x8m81_0/xb[0] xdec64_3v256x8m81_0/xa[7]
+ xdec64_3v256x8m81_0/xa[6] xdec64_3v256x8m81_0/xa[5] xdec64_3v256x8m81_0/xa[4] xdec64_3v256x8m81_0/xa[2]
+ A[0] xdec64_3v256x8m81_0/xb[1] control_3v256x8_3v256x8m81_0/xc[3] xdec64_3v256x8m81_0/xc[1]
+ control_3v256x8_3v256x8m81_0/xc[2] xdec64_3v256x8m81_0/xa[1] VSS A[7] CLK A[2] A[1]
+ A[6] A[3] A[4] A[5] VSS rcol4_256_3v256x8m81_0/GWE GWEN lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[1]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[2] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[4]
+ xdec64_3v256x8m81_0/xa[3] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[5]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[6] xdec64_3v256x8m81_0/xa[0]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[7] CEN control_3v256x8_3v256x8m81_0/xc[0]
+ xdec64_3v256x8m81_0/men VDD VSS VDD control_3v256x8_3v256x8m81
Xxdec64_3v256x8m81_0 xdec64_3v256x8m81_0/DRWL xdec64_3v256x8m81_0/DLWL xdec64_3v256x8m81_0/LWL[20]
+ xdec64_3v256x8m81_0/LWL[21] xdec64_3v256x8m81_0/LWL[22] xdec64_3v256x8m81_0/LWL[27]
+ xdec64_3v256x8m81_0/LWL[13] xdec64_3v256x8m81_0/LWL[14] xdec64_3v256x8m81_0/LWL[16]
+ xdec64_3v256x8m81_0/LWL[3] xdec64_3v256x8m81_0/LWL[2] xdec64_3v256x8m81_0/LWL[1]
+ xdec64_3v256x8m81_0/LWL[0] xdec64_3v256x8m81_0/LWL[8] xdec64_3v256x8m81_0/LWL[9]
+ xdec64_3v256x8m81_0/LWL[7] xdec64_3v256x8m81_0/LWL[30] xdec64_3v256x8m81_0/RWL[31]
+ xdec64_3v256x8m81_0/RWL[30] xdec64_3v256x8m81_0/RWL[29] xdec64_3v256x8m81_0/RWL[22]
+ xdec64_3v256x8m81_0/RWL[4] xdec64_3v256x8m81_0/RWL[2] xdec64_3v256x8m81_0/RWL[0]
+ xdec64_3v256x8m81_0/RWL[1] xdec64_3v256x8m81_0/RWL[3] xdec64_3v256x8m81_0/RWL[7]
+ xdec64_3v256x8m81_0/RWL[9] xdec64_3v256x8m81_0/RWL[11] xdec64_3v256x8m81_0/RWL[14]
+ xdec64_3v256x8m81_0/RWL[15] xdec64_3v256x8m81_0/RWL[16] xdec64_3v256x8m81_0/RWL[17]
+ xdec64_3v256x8m81_0/RWL[18] xdec64_3v256x8m81_0/RWL[19] xdec64_3v256x8m81_0/RWL[20]
+ xdec64_3v256x8m81_0/xb[0] xdec64_3v256x8m81_0/xb[1] xdec64_3v256x8m81_0/xb[2] xdec64_3v256x8m81_0/xb[3]
+ xdec64_3v256x8m81_0/xa[7] xdec64_3v256x8m81_0/xa[6] xdec64_3v256x8m81_0/xa[5] xdec64_3v256x8m81_0/xa[4]
+ xdec64_3v256x8m81_0/xa[0] xdec64_3v256x8m81_0/men xdec64_3v256x8m81_0/xa[3] xdec64_3v256x8m81_0/xa[2]
+ xdec64_3v256x8m81_0/xa[1] xdec64_3v256x8m81_0/xc[1] xdec64_3v256x8m81_0/RWL[21]
+ xdec64_3v256x8m81_0/LWL[25] xdec64_3v256x8m81_0/LWL[28] xdec64_3v256x8m81_0/LWL[26]
+ xdec64_3v256x8m81_0/LWL[11] xdec64_3v256x8m81_0/LWL[12] xdec64_3v256x8m81_0/LWL[24]
+ xdec64_3v256x8m81_0/RWL[27] xdec64_3v256x8m81_0/LWL[23] xdec64_3v256x8m81_0/LWL[10]
+ xdec64_3v256x8m81_0/LWL[31] xdec64_3v256x8m81_0/LWL[19] xdec64_3v256x8m81_0/RWL[12]
+ xdec64_3v256x8m81_0/LWL[17] xdec64_3v256x8m81_0/RWL[28] xdec64_3v256x8m81_0/RWL[25]
+ VDD xdec64_3v256x8m81_0/RWL[10] xdec64_3v256x8m81_0/LWL[29] xdec64_3v256x8m81_0/RWL[5]
+ xdec64_3v256x8m81_0/RWL[26] VSS xdec64_3v256x8m81_0/LWL[5] xdec64_3v256x8m81_0/LWL[6]
+ xdec64_3v256x8m81_0/RWL[13] xdec64_3v256x8m81_0/LWL[18] xdec64_3v256x8m81_0/RWL[24]
+ xdec64_3v256x8m81_0/RWL[8] xdec64_3v256x8m81_0/LWL[4] xdec64_3v256x8m81_0/LWL[15]
+ VDD xdec64_3v256x8m81_0/RWL[23] xdec64_3v256x8m81_0/RWL[6] xdec64_3v256x8m81
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__mux2_4 VDD VNW VPW VSS S B A Y
X0 a_744_440# S a_464_68# VNW pfet_03v3 ad=0.1932p pd=1.66u as=0.3588p ps=1.9u w=1.38u l=0.28u
X1 VDD A a_744_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.1932p ps=1.66u w=1.38u l=0.28u
X2 VDD a_464_68# Y VNW pfet_03v3 ad=0.828p pd=3.96u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 a_332_440# B VDD VNW pfet_03v3 ad=0.6762p pd=2.36u as=0.3588p ps=1.9u w=1.38u l=0.28u
X4 a_464_68# S a_332_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.19p ps=1.38u w=1u l=0.28u
X5 VSS S a_28_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 Y a_464_68# VDD VNW pfet_03v3 ad=0.3726p pd=1.92u as=0.3588p ps=1.9u w=1.38u l=0.28u
X7 Y a_464_68# VSS VPW nfet_03v3 ad=0.27p pd=1.54u as=0.26p ps=1.52u w=1u l=0.28u
X8 VSS a_464_68# Y VPW nfet_03v3 ad=0.6p pd=3.2u as=0.26p ps=1.52u w=1u l=0.28u
X9 VSS A a_624_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=1.88u w=1u l=0.28u
X10 VDD a_464_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3726p ps=1.92u w=1.38u l=0.28u
X11 Y a_464_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 Y a_464_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X13 VSS a_464_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.27p ps=1.54u w=1u l=0.28u
X14 a_464_68# a_28_68# a_332_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6762p ps=2.36u w=1.38u l=0.28u
X15 VDD S a_28_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X16 a_624_68# a_28_68# a_464_68# VPW nfet_03v3 ad=0.44p pd=1.88u as=0.26p ps=1.52u w=1u l=0.28u
X17 a_332_68# B VSS VPW nfet_03v3 ad=0.19p pd=1.38u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__fillcap_4 VDD VNW VPW VSS
X0 a_126_408# a_28_500# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.49p ps=2.98u w=1u l=1.03u
X1 VDD a_126_408# a_28_500# VNW pfet_03v3 ad=0.4752p pd=3.04u as=0.5292p ps=3.14u w=1.08u l=1.03u
.ends

.subckt ocd_mux_array S A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[7] B[6] B[5] B[4]
+ B[3] B[2] B[1] B[0] Y[7] Y[3] Y[5] Y[1] Y[6] vdd Y[4] Y[0] vss Y[2]
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_8 vdd vdd vss vss S B[6] A[6] Y[6] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_9 vdd vdd vss vss S B[7] A[7] Y[7] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__fillcap_4_2 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__fillcap_4
Xgf180mcu_as_sc_mcu7t3v3__fillcap_4_3 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__fillcap_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_10 vdd vdd vss vss S B[3] A[3] Y[3] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_11 vdd vdd vss vss S B[4] A[4] Y[4] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_12 vdd vdd vss vss S B[5] A[5] Y[5] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_13 vdd vdd vss vss S B[0] A[0] Y[0] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_14 vdd vdd vss vss S B[1] A[1] Y[1] gf180mcu_as_sc_mcu7t3v3__mux2_4
Xgf180mcu_as_sc_mcu7t3v3__mux2_4_15 vdd vdd vss vss S B[2] A[2] Y[2] gf180mcu_as_sc_mcu7t3v3__mux2_4
.ends

.subckt POLY_SUB_FILL_1 a_597_223# a_685_131#
X0 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
X1 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
.ends

.subckt GF_NI_FILL10_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[14] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[15] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0 DVSS DVDD VDD VSS
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1
.ends

.subckt gf180mcu_ocd_io__fill10 VDD VSS DVDD DVSS
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0
.ends

.subckt POLY_SUB_FILL a_1165_n91# a_1077_1#
X0 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
X1 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
.ends

.subckt GF_NI_FILL5_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_0[0] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[1] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[2] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[3] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[4] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[5] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[6] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[7] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[8] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[9] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[10] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[11] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[12] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[13] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[14] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[15] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[16] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[17] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[18] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[19] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[20] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[21] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[22] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[23] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[24] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[25] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[26] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[27] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[28] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[29] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[30] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[31] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[32] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[33] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[34] VDD VSS POLY_SUB_FILL
.ends

.subckt GF_NI_FILL5_0 DVSS DVDD VDD VSS
XGF_NI_FILL5_1_0 VSS VDD DVSS DVDD GF_NI_FILL5_1
.ends

.subckt gf180mcu_ocd_io__fill5 VDD VSS DVDD DVSS
XGF_NI_FILL5_0_0 DVSS DVDD VDD VSS GF_NI_FILL5_0
.ends

.subckt lv_nand a_16960_50788# w_16870_51136# a_17113_51095# a_17024_51222# a_17252_51095#
X0 a_17204_50930# a_17113_51095# a_16960_50788# a_16960_50788# nfet_03v3 ad=0.114p pd=0.98u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_17024_51222# a_17252_51095# a_17204_50930# a_16960_50788# nfet_03v3 ad=0.264p pd=2.08u as=0.114p ps=0.98u w=0.6u l=0.28u
X2 w_16870_51136# a_17113_51095# a_17024_51222# w_16870_51136# pfet_03v3 ad=0.333p pd=1.755u as=0.534p ps=3.29u w=1.2u l=0.28u
X3 a_17024_51222# a_17252_51095# w_16870_51136# w_16870_51136# pfet_03v3 ad=0.528p pd=3.28u as=0.333p ps=1.755u w=1.2u l=0.28u
.ends

.subckt pmos_6p0_esd_40 w_0_12# a_278_44# a_974_132# a_222_132#
X0 a_974_132# a_278_44# a_222_132# w_0_12# pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.2p ps=80.56u w=40u l=0.7u
.ends

.subckt comp018green_out_drv_pleg_4T_Y pmos_6p0_esd_40_0/w_0_12# pmos_6p0_esd_40_0/a_278_44#
+ pmos_6p0_esd_40_0/a_974_132# pmos_6p0_esd_40_0/a_222_132#
Xpmos_6p0_esd_40_0 pmos_6p0_esd_40_0/w_0_12# pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_0/a_974_132#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40
.ends

.subckt comp018green_out_drv_pleg_4T_X pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_1/w_0_12#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40_1/a_974_132# pmos_6p0_esd_40_1/a_278_44#
+ pmos_6p0_esd_40_1/a_222_132#
Xpmos_6p0_esd_40_0 pmos_6p0_esd_40_1/w_0_12# pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_1/a_974_132#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40
Xpmos_6p0_esd_40_1 pmos_6p0_esd_40_1/w_0_12# pmos_6p0_esd_40_1/a_278_44# pmos_6p0_esd_40_1/a_974_132#
+ pmos_6p0_esd_40_1/a_222_132# pmos_6p0_esd_40
.ends

.subckt comp018green_out_paddrv_4T_PMOS_GROUP PMOS_4T_metal_stack_4/m1_340_0# a_2360_2800#
+ PMOS_4T_metal_stack_5/m1_340_0# a_4511_2800# PMOS_4T_metal_stack_5/m1_n44_0# PMOS_4T_metal_stack_1/m1_n44_0#
+ PMOS_4T_metal_stack_1/m1_340_0# PMOS_4T_metal_stack_2/m1_n44_0# a_9428_2800# a_7662_2800#
+ a_11201_2800# a_9815_2800# PMOS_4T_metal_stack_6/m1_340_0# PMOS_4T_metal_stack_2/m1_340_0#
+ PMOS_4T_metal_stack_3/m1_n44_0# a_6280_2800# a_2746_2800# a_974_2800# a_8049_2800#
+ a_5892_2800# PMOS_4T_metal_stack_3/m1_340_0# a_4120_2800# PMOS_4T_metal_stack_4/m1_n44_0#
+ w_n5_111#
Xcomp018green_out_drv_pleg_4T_Y_0 w_n5_111# a_4120_2800# PMOS_4T_metal_stack_1/m1_340_0#
+ PMOS_4T_metal_stack_2/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_1 w_n5_111# a_9428_2800# PMOS_4T_metal_stack_4/m1_340_0#
+ PMOS_4T_metal_stack_5/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_2 w_n5_111# a_2746_2800# PMOS_4T_metal_stack_1/m1_340_0#
+ PMOS_4T_metal_stack_1/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_3 w_n5_111# a_8049_2800# PMOS_4T_metal_stack_4/m1_340_0#
+ PMOS_4T_metal_stack_4/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_X_0 a_4511_2800# w_n5_111# PMOS_4T_metal_stack_2/m1_n44_0#
+ PMOS_4T_metal_stack_2/m1_340_0# a_5892_2800# PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_1 a_9815_2800# w_n5_111# PMOS_4T_metal_stack_5/m1_n44_0#
+ PMOS_4T_metal_stack_5/m1_340_0# a_11201_2800# w_n5_111# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_2 a_7662_2800# w_n5_111# PMOS_4T_metal_stack_4/m1_n44_0#
+ PMOS_4T_metal_stack_3/m1_340_0# a_6280_2800# PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_3 a_2360_2800# w_n5_111# PMOS_4T_metal_stack_1/m1_n44_0#
+ PMOS_4T_metal_stack_6/m1_340_0# a_974_2800# w_n5_111# comp018green_out_drv_pleg_4T_X
.ends

.subckt comp018green_out_drv_nleg_4T a_206_444# a_2080_444# a_2366_532# a_48_532#
+ a_436_532# VSUBS
X0 a_436_532# a_206_444# a_48_532# VSUBS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.64p ps=76.56u w=38u l=1.15u
X1 a_2366_532# a_2080_444# a_436_532# VSUBS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.64p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
.ends

.subckt comp018green_out_paddrv_4T_NMOS_GROUP GR_NMOS_4T_0/w_n1730_n583# a_7847_1028#
+ a_7373_1028# a_803_1028# nmos_4T_metal_stack_1/m1_n44_400# nmos_4T_metal_stack_2/m1_n44_400#
+ nmos_4T_metal_stack_3/m1_n44_400# nmos_4T_metal_stack_3/m1_430_401# a_2677_1028#
+ nmos_4T_metal_stack_1/m1_430_401# a_9721_1028# nmos_4T_metal_stack_2/m1_430_401#
+ nmos_4T_metal_stack_0/m1_n44_400# nmos_4T_metal_stack_4/m1_430_401# a_5499_1028#
+ a_3151_1028# VSUBS a_5025_1028# nmos_4T_metal_stack_4/m1_n44_400#
Xcomp018green_out_drv_nleg_4T_0 a_7847_1028# a_9721_1028# nmos_4T_metal_stack_0/m1_n44_400#
+ nmos_4T_metal_stack_3/m1_n44_400# nmos_4T_metal_stack_3/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_1 a_5499_1028# a_7373_1028# nmos_4T_metal_stack_3/m1_n44_400#
+ nmos_4T_metal_stack_2/m1_n44_400# nmos_4T_metal_stack_2/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_2 a_3151_1028# a_5025_1028# nmos_4T_metal_stack_2/m1_n44_400#
+ nmos_4T_metal_stack_1/m1_n44_400# nmos_4T_metal_stack_1/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_3 a_803_1028# a_2677_1028# nmos_4T_metal_stack_1/m1_n44_400#
+ nmos_4T_metal_stack_4/m1_n44_400# nmos_4T_metal_stack_4/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
.ends

.subckt comp018green_out_paddrv_16T comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800#
+ m1_12305_8954# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800# m1_n360_8434# m1_1026_8954#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0# m1_12305_9280#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400# m1_12305_9120#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800# m1_1026_9280# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ m1_1026_9120# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m1_12305_9446# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# m2_1697_23319#
+ m1_1026_9446# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
Xcomp018green_out_paddrv_4T_PMOS_GROUP_0 m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0# m2_1697_23319#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800# m2_1697_23319# m2_1697_23319#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111# comp018green_out_paddrv_4T_PMOS_GROUP
Xcomp018green_out_paddrv_4T_NMOS_GROUP_0 m1_n360_8434# m1_12305_9120# m1_12305_9280#
+ m1_1026_8954# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ m2_1697_23319# m1_1026_9120# m2_1697_23319# m1_12305_8954# m2_1697_23319# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m2_1697_23319# m1_12305_9446# m1_1026_9280# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m1_1026_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS comp018green_out_paddrv_4T_NMOS_GROUP
.ends

.subckt tie_poly_res a_n2051_55943# a_n2051_55061# a_n2331_55943# w_n2756_54700#
X0 a_n2051_55943# a_n2051_55061# w_n2756_54700# ppolyf_u r_width=0.8u r_length=3.9u
X1 a_n2331_55943# w_n2756_54700# w_n2756_54700# ppolyf_u r_width=0.8u r_length=3.9u
.ends

.subckt lvlshift_up a_18491_55181# a_18216_53410# a_18479_54386# a_18481_54667# w_18130_54691#
X0 w_18130_54691# a_18491_55181# a_18403_53764# w_18130_54691# pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X1 a_18491_55181# a_18403_53764# w_18130_54691# w_18130_54691# pfet_06v0 ad=0.675p pd=3.9u as=0.39p ps=2.02u w=1.5u l=0.7u
X2 a_18216_53410# a_18479_54386# a_18403_53764# a_18216_53410# nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X3 a_18491_55181# a_18481_54667# a_18216_53410# a_18216_53410# nfet_06v0 ad=0.675p pd=3.9u as=0.39p ps=2.02u w=1.5u l=0.7u
.ends

.subckt comp018green_sigbuf_1 Z DVSS DVDD ZB lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1605_310# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 DVSS Z ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 Z a_1605_310# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X2 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X4 ZB Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X5 DVDD a_1605_310# Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X6 Z a_1605_310# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X7 DVSS a_1605_310# Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
.ends

.subckt comp018green_out_predrv SL SLB NDRIVE_X ENB DVSS A DVDD NDRIVE_Y PDRIVE_Y
+ PDRIVE_X EN
X0 a_1395_3267# ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X1 DVDD a_1395_3267# PDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X2 NDRIVE_X a_335_226# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X3 a_335_226# EN a_1395_3267# DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X4 NDRIVE_Y SL NDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X5 DVSS a_335_226# NDRIVE_X DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X6 a_335_226# A DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X7 DVDD a_335_226# NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X8 PDRIVE_X a_1395_3267# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X9 PDRIVE_X DVDD PDRIVE_Y DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X10 PDRIVE_Y SLB PDRIVE_X DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X11 NDRIVE_Y a_335_226# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X12 PDRIVE_X SLB PDRIVE_Y DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X13 NDRIVE_Y a_335_226# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X14 a_335_226# ENB a_1395_3267# DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X15 DVDD EN a_335_226# DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X16 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X17 DVSS A a_1395_3267# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X18 DVSS a_335_226# NDRIVE_Y DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X19 DVDD a_1395_3267# PDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X20 PDRIVE_Y a_1395_3267# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X21 PDRIVE_Y a_1395_3267# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X22 DVSS a_1395_3267# PDRIVE_Y DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X23 NDRIVE_X SL NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
.ends

.subckt comp018green_out_sigbuf_a AB DVSS DVDD lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1697_1072# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 AB a_1825_270# DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X1 AB a_1825_270# DVDD DVDD pfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X2 DVSS a_1697_1072# a_1825_270# DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X3 DVDD a_1697_1072# a_1825_270# DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
.ends

.subckt comp018green_out_sigbuf_oe ENB DVDD DVSS EN lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1783_1072# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 DVDD a_1783_1072# EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X1 DVSS a_1783_1072# EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X2 ENB EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X3 ENB EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt lv_inv w_15980_51147# a_16280_50941# a_16119_51106# a_16066_50799#
X0 a_16280_50941# a_16119_51106# a_16066_50799# a_16066_50799# nfet_03v3 ad=0.264p pd=2.08u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_16280_50941# a_16119_51106# w_15980_51147# w_15980_51147# pfet_03v3 ad=0.528p pd=3.28u as=0.558p ps=3.33u w=1.2u l=0.28u
.ends

.subckt comp018green_in_pupd A DVDD DVSS PU_B PD w_n83_53# a_506_484# a_6234_n7404#
X0 DVSS PD a_6278_n7492# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X1 a_404_1044# a_7646_1324# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X2 a_404_2164# a_6278_n7492# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X3 DVDD a_6234_n7404# a_6278_n7492# DVDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X4 a_404_484# a_7646_764# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X5 a_404_1044# a_7646_764# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X6 a_404_2164# a_7646_1884# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X7 a_404_484# A w_n83_53# ppolyf_u r_width=0.8u r_length=23u
X8 a_404_1604# a_7646_1884# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X9 a_404_1604# a_7646_1324# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
.ends

.subckt lv_passgate a_15637_45872# a_15397_45912# w_15280_46078# a_15366_45730# a_15492_45872#
+ a_15396_46108#
X0 a_15637_45872# a_15397_45912# a_15492_45872# a_15366_45730# nfet_03v3 ad=0.264p pd=2.08u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_15637_45872# a_15396_46108# a_15492_45872# w_15280_46078# pfet_03v3 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.28u
.ends

.subckt comp018green_in_logic_pupd m1_1586_653# m1_1573_n494# m1_1324_578# m1_1842_n2708#
+ m1_1316_n577# a_1638_n204# w_1648_203# m1_1455_n1573#
Xlv_nand_4 a_1638_n204# w_1648_203# m1_1842_n2708# m1_1921_n496# m1_1909_n1494# lv_nand
Xlv_inv_0 w_1648_203# m1_1573_n494# m1_1921_n496# a_1638_n204# lv_inv
Xlv_inv_1 w_1648_203# m1_1586_653# m1_1910_652# a_1638_n204# lv_inv
Xlv_inv_2 w_1648_203# m1_1455_n1773# m1_1455_n1573# a_1638_n204# lv_inv
Xlv_passgate_0 m1_1909_n1494# m1_1455_n1573# w_1648_203# a_1638_n204# m1_1580_n1918#
+ m1_1455_n1773# lv_passgate
Xlv_inv_3 w_1648_203# m1_1580_n1918# m1_1842_n2708# a_1638_n204# lv_inv
Xlv_passgate_1 m1_1909_n1494# m1_1455_n1773# w_1648_203# a_1638_n204# m1_1842_n2708#
+ m1_1455_n1573# lv_passgate
Xlv_inv_5 w_1648_203# m1_1324_578# m1_1586_653# a_1638_n204# lv_inv
Xlv_inv_7 w_1648_203# m1_1316_n577# m1_1573_n494# a_1638_n204# lv_inv
Xlv_nand_0 a_1638_n204# w_1648_203# m1_1455_n1573# m1_1910_652# m1_1909_n1494# lv_nand
.ends

.subckt comp018green_sigbuf Z DVSS DVDD ZB INB IN
Xlvlshift_up_0 a_1561_310# DVSS IN INB DVDD lvlshift_up
X0 ZB Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 DVSS Z ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X2 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVSS a_1561_310# Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X4 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X5 Z a_1561_310# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X6 Z a_1561_310# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X7 DVDD a_1561_310# Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt comp018green_in_drv A VDD VSS Z a_2771_580# a_1167_270# w_2679_1281# a_923_1522#
+ a_3067_747#
X0 VSS A a_n180_263# VSS nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X1 a_n180_263# A VSS VSS nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X2 Z a_n180_263# a_1167_270# VSS nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
X3 a_1167_270# a_n180_263# Z VSS nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X4 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X5 a_923_1522# a_n180_263# Z VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X6 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X7 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.644p ps=3.72u w=1.4u l=0.28u
X8 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.276p ps=2.12u w=0.6u l=0.28u
X9 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X10 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X11 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.276p pd=2.12u as=0.162p ps=1.14u w=0.6u l=0.28u
X12 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X13 Z a_n180_263# a_923_1522# VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X14 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.644p pd=3.72u as=0.378p ps=1.94u w=1.4u l=0.28u
X15 a_n180_263# A VDD VDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X16 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X17 a_923_1522# a_n180_263# Z VDD pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
X18 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X19 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X20 Z a_n180_263# a_923_1522# VDD pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
.ends

.subckt comp018green_in_cms_smt IE CS DVDD A DVSS Z a_5355_608# m2_5364_1052#
X0 a_1887_280# IE DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X1 a_3115_338# a_1082_620# a_5355_608# DVSS nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X2 a_1082_620# a_599_280# Z DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X3 DVSS CS a_599_280# DVSS nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X4 DVSS a_1809_1797# a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X5 DVSS IE a_1887_280# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X6 Z CS a_1809_1797# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X7 Z IE DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X8 Z a_599_280# a_1809_1797# DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X9 a_1887_280# A a_3115_338# DVSS nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
X10 DVDD CS a_1809_1797# DVDD pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X11 a_3115_338# A a_1887_280# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X12 Z A a_3227_1730# DVDD pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X13 a_3227_1730# A Z DVDD pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X14 DVSS a_599_280# a_1082_620# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X15 a_1887_280# A a_3115_338# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X16 DVDD A a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X17 a_1887_280# IE DVSS DVSS nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X18 Z A a_3115_338# DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X19 a_599_280# CS DVDD DVDD pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X20 Z IE DVDD DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X21 a_3115_338# A Z DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X22 DVDD IE Z DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X23 a_3115_338# A a_1887_280# DVSS nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X24 a_1082_620# CS Z DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X25 a_3227_1730# A DVDD DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X26 a_3115_338# A Z DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X27 a_3227_1730# a_1809_1797# DVSS DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X28 a_599_280# CS DVSS DVSS nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X29 DVDD CS a_599_280# DVDD pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X30 a_1887_280# IE DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
X31 Z A a_3115_338# DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X32 a_1809_1797# CS DVDD DVDD pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X33 DVSS IE a_1887_280# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
.ends

.subckt comp018green_inpath_cms_smt PAD CS PU comp018green_in_cms_smt_0/a_5355_608#
+ a_1390_1224# comp018green_in_logic_pupd_0/w_1648_203# comp018green_in_pupd_0/w_n83_53#
+ comp018green_in_pupd_0/A m3_9619_4882# m3_9619_3696# comp018green_in_pupd_0/DVSS
+ comp018green_in_pupd_0/DVDD comp018green_in_drv_0/VDD comp018green_in_drv_0/VSS
+ m1_12910_4326# VSUBS m1_10570_5335# comp018green_in_pupd_0/a_506_484# a_1390_2124#
+ w_n13_970# comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
Xlv_inv_14 w_n13_970# comp018green_sigbuf_1/IN a_1390_1224# VSUBS lv_inv
Xlv_inv_15 w_n13_970# comp018green_sigbuf_1/INB comp018green_sigbuf_1/IN VSUBS lv_inv
Xcomp018green_in_pupd_0 comp018green_in_pupd_0/A comp018green_in_pupd_0/DVDD comp018green_in_pupd_0/DVSS
+ comp018green_in_pupd_0/PU_B comp018green_sigbuf_0/ZB comp018green_in_pupd_0/w_n83_53#
+ comp018green_in_pupd_0/a_506_484# comp018green_sigbuf_2/Z comp018green_in_pupd
Xcomp018green_in_logic_pupd_0 comp018green_sigbuf_0/IN comp018green_sigbuf_2/IN comp018green_sigbuf_0/INB
+ PU comp018green_sigbuf_2/INB VSUBS comp018green_in_logic_pupd_0/w_1648_203# a_1390_2124#
+ comp018green_in_logic_pupd
Xcomp018green_sigbuf_0 comp018green_sigbuf_0/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_0/ZB comp018green_sigbuf_0/INB comp018green_sigbuf_0/IN comp018green_sigbuf
Xlv_inv_18 w_n13_970# comp018green_sigbuf_3/IN CS VSUBS lv_inv
Xlv_inv_19 w_n13_970# comp018green_sigbuf_3/INB comp018green_sigbuf_3/IN VSUBS lv_inv
Xcomp018green_sigbuf_1 comp018green_sigbuf_1/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_1/ZB comp018green_sigbuf_1/INB comp018green_sigbuf_1/IN comp018green_sigbuf
Xcomp018green_sigbuf_2 comp018green_sigbuf_2/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_2/ZB comp018green_sigbuf_2/INB comp018green_sigbuf_2/IN comp018green_sigbuf
Xcomp018green_sigbuf_3 comp018green_sigbuf_3/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_3/ZB comp018green_sigbuf_3/INB comp018green_sigbuf_3/IN comp018green_sigbuf
Xcomp018green_in_drv_0 comp018green_in_drv_0/A comp018green_in_drv_0/VDD comp018green_in_drv_0/VSS
+ comp018green_in_drv_0/Z VSUBS VSUBS m1_10570_5335# m1_10570_5335# m1_12910_4326#
+ comp018green_in_drv
Xcomp018green_in_cms_smt_0 comp018green_sigbuf_1/Z comp018green_sigbuf_3/Z comp018green_in_drv_0/VDD
+ PAD comp018green_in_drv_0/VSS comp018green_in_drv_0/A comp018green_in_cms_smt_0/a_5355_608#
+ PAD comp018green_in_cms_smt
D0 CS w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D1 a_1390_1224# w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D2 PU w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D3 a_1390_2124# w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
.ends

.subckt comp018green_esd_cdm IP_IN PAD DVDD DVSS w_n86_n86# w_454_3720#
X0 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
D0 DVSS IP_IN diode_nd2ps_06v0 pj=42u area=20p
D1 IP_IN w_454_3720# diode_pd2nw_06v0 pj=42u area=20p
D2 DVSS IP_IN diode_nd2ps_06v0 pj=42u area=20p
X1 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
X2 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
X3 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
D3 IP_IN w_454_3720# diode_pd2nw_06v0 pj=42u area=20p
.ends

.subckt GF_NI_IN_C_BASE PD PU Y ndrive_y_<0> ndrive_x_<0> ndrive_x_<1> ndrive_Y_<1>
+ ndrive_x_<2> ndrive_y_<2> ndrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_y_<0> pdrive_y_<1>
+ pdrive_x_<1> pdrive_x_<2> pdrive_y_<2> pdrive_y_<3> pdrive_x_<3> m3_1771_39126#
+ w_11000_43887# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ m2_1886_52816# comp018green_inpath_cms_smt_0/m3_9619_4882# w_873_53312# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_esd_cdm_0/w_454_3720# m3_10025_37504# PAD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ a_12390_41548# m1_3608_46684# comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ tie_poly_res_0/VSUBS comp018green_sigbuf_1_0/DVSS comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_sigbuf_1_0/DVDD comp018green_inpath_cms_smt_0/m1_10570_5335# comp018green_inpath_cms_smt_0/VSUBS
+ w_11042_41027# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_predrv_3/DVDD w_13720_39292# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
Xlv_nand_2 tie_poly_res_0/VSUBS w_13720_39292# comp018green_inpath_cms_smt_0/CS m1_5236_36986#
+ w_13720_39292# lv_nand
Xlv_nand_3 tie_poly_res_0/VSUBS w_13720_39292# comp018green_inpath_cms_smt_0/CS m1_4812_38523#
+ comp018green_inpath_cms_smt_0/CS lv_nand
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ pdrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> comp018green_out_predrv_3/DVDD
+ ndrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ ndrive_y_<2> pdrive_y_<2> pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ ndrive_y_<0> pdrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ ndrive_x_<2> pdrive_x_<1> PAD ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_out_paddrv_16T
Xtie_poly_res_0 comp018green_inpath_cms_smt_0/CS comp018green_inpath_cms_smt_0/VSUBS
+ m1_1554_56149# w_873_53312# tie_poly_res
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/DVSS comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/ZB m1_9774_36986# m1_9537_37107# comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<0> pdrive_y_<0> pdrive_x_<0> comp018green_out_predrv_0/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD m1_9174_38525# m1_9257_38818# comp018green_out_sigbuf_a
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<2> pdrive_y_<2> pdrive_x_<2> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<3> pdrive_y_<3> pdrive_x_<3> comp018green_out_predrv_1/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_0/EN m1_1182_38534# m1_1187_38806#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<1> pdrive_y_<1> pdrive_x_<1> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/CS
+ PU comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD m1_1554_56149# w_11000_43887#
+ m1_3608_46684# comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/m3_9619_4882#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
+ Y comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/m1_10570_5335#
+ comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484# PD w_873_53312#
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_1/EN m1_5236_36986# m1_5084_37107#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_sigbuf_oe_1 comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/EN m1_4812_38523# m1_4626_36747#
+ comp018green_out_sigbuf_oe
Xlv_inv_0 w_13720_39292# m1_1187_38806# m1_1182_38534# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_1 w_13720_39292# m1_9257_38818# m1_9174_38525# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_2 w_13720_39292# m1_9537_37107# m1_9774_36986# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_3 w_13720_39292# m1_4626_36747# m1_4812_38523# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_4 w_13720_39292# m1_9774_36986# comp018green_inpath_cms_smt_0/CS tie_poly_res_0/VSUBS
+ lv_inv
Xlv_inv_6 w_13720_39292# m1_5084_37107# m1_5236_36986# tie_poly_res_0/VSUBS lv_inv
Xcomp018green_esd_cdm_0 comp018green_esd_cdm_0/IP_IN PAD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm
Xlv_nand_0 tie_poly_res_0/VSUBS w_13720_39292# comp018green_inpath_cms_smt_0/CS m1_9174_38525#
+ comp018green_inpath_cms_smt_0/CS lv_nand
Xlv_nand_1 tie_poly_res_0/VSUBS w_13720_39292# comp018green_inpath_cms_smt_0/CS m1_1182_38534#
+ comp018green_inpath_cms_smt_0/CS lv_nand
X0 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X1 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X2 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X4 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X5 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X6 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X7 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X8 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X9 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
D0 comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS diode_pd2nw_03v3 pj=1.92u area=0.2304p
D1 comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS diode_pd2nw_03v3 pj=1.92u area=0.2304p
D2 comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS diode_pd2nw_03v3 pj=1.92u area=0.2304p
D3 comp018green_inpath_cms_smt_0/VSUBS w_11000_43887# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D4 comp018green_inpath_cms_smt_0/CS w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
D5 comp018green_inpath_cms_smt_0/CS w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
X10 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
D6 comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS diode_pd2nw_03v3 pj=1.92u area=0.2304p
D7 comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS diode_pd2nw_03v3 pj=1.92u area=0.2304p
X11 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt gf180mcu_ocd_io__in_c DVDD PD PU VDD Y PAD DVSS VSS
XGF_NI_IN_C_BASE_0 PD PU Y GF_NI_IN_C_BASE_0/ndrive_y_<0> GF_NI_IN_C_BASE_0/ndrive_x_<0>
+ GF_NI_IN_C_BASE_0/ndrive_x_<1> GF_NI_IN_C_BASE_0/ndrive_Y_<1> GF_NI_IN_C_BASE_0/ndrive_x_<2>
+ GF_NI_IN_C_BASE_0/ndrive_y_<2> GF_NI_IN_C_BASE_0/ndrive_x_<3> GF_NI_IN_C_BASE_0/ndrive_Y_<3>
+ GF_NI_IN_C_BASE_0/pdrive_x_<0> GF_NI_IN_C_BASE_0/pdrive_y_<0> GF_NI_IN_C_BASE_0/pdrive_y_<1>
+ GF_NI_IN_C_BASE_0/pdrive_x_<1> GF_NI_IN_C_BASE_0/pdrive_x_<2> GF_NI_IN_C_BASE_0/pdrive_y_<2>
+ GF_NI_IN_C_BASE_0/pdrive_y_<3> GF_NI_IN_C_BASE_0/pdrive_x_<3> VDD VDD DVDD DVDD
+ DVSS VDD VDD DVSS VSS DVSS DVSS DVDD DVDD DVDD VSS PAD DVDD DVDD DVDD DVDD DVDD
+ DVDD VSS DVSS DVSS DVDD DVDD VDD VSS VDD DVSS DVDD VDD DVSS GF_NI_IN_C_BASE
.ends

.subckt GF_NI_BI_T_BASE PD IE SL A OE CS PU PDRV0 PDRV1 Y ndrive_y_<0> ndrive_x_<0>
+ ndrive_x_<1> ndrive_Y_<1> ndrive_x_<2> ndrive_y_<2> ndrive_x_<3> ndrive_Y_<3> pdrive_x_<0>
+ pdrive_y_<0> pdrive_y_<1> pdrive_x_<1> pdrive_x_<2> pdrive_y_<2> pdrive_y_<3> pdrive_x_<3>
+ m3_1771_39126# w_11000_43887# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_inpath_cms_smt_0/m3_9619_4882# w_835_53274# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_esd_cdm_0/w_454_3720# m3_10025_37504# PAD comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ a_12390_41548# m1_3608_46684# comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_sigbuf_1_0/VSUBS comp018green_esd_cdm_0/IP_IN comp018green_sigbuf_1_0/DVSS
+ comp018green_esd_cdm_0/DVSS comp018green_sigbuf_1_0/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ a_882_55933# comp018green_inpath_cms_smt_0/m1_10570_5335# comp018green_inpath_cms_smt_0/VSUBS
+ w_11042_41027# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_predrv_3/DVDD w_13720_39292# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
Xlv_nand_2 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_5236_36986# w_13720_39292#
+ lv_nand
Xlv_nand_3 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_4812_38523# PDRV1 lv_nand
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ pdrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> comp018green_out_predrv_3/DVDD
+ ndrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ ndrive_y_<2> pdrive_y_<2> pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ ndrive_y_<0> pdrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ ndrive_x_<2> pdrive_x_<1> PAD ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_out_paddrv_16T
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/DVSS comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/ZB m1_9774_36986# m1_9537_37107# comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<0> pdrive_y_<0> pdrive_x_<0> comp018green_out_predrv_0/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD m1_9178_38525# m1_9257_38818# comp018green_out_sigbuf_a
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<2> pdrive_y_<2> pdrive_x_<2> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<3> pdrive_y_<3> pdrive_x_<3> comp018green_out_predrv_1/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_0/EN m1_1184_38534# m1_1189_38806#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<1> pdrive_y_<1> pdrive_x_<1> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN CS PU comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ IE w_11000_43887# m1_3608_46684# comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/m3_9619_4882#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
+ Y comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/m1_10570_5335#
+ comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484# PD w_835_53274#
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_1/EN m1_5236_36986# m1_5084_37107#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_sigbuf_oe_1 comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/EN m1_4812_38523# m1_4626_36747#
+ comp018green_out_sigbuf_oe
Xlv_inv_0 w_13720_39292# m1_1189_38806# m1_1184_38534# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_1 w_13720_39292# m1_9257_38818# m1_9178_38525# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_2 w_13720_39292# m1_9537_37107# m1_9774_36986# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_3 w_13720_39292# m1_4626_36747# m1_4812_38523# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_4 w_13720_39292# m1_9774_36986# SL comp018green_sigbuf_1_0/VSUBS lv_inv
Xlv_inv_6 w_13720_39292# m1_5084_37107# m1_5236_36986# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xcomp018green_esd_cdm_0 comp018green_esd_cdm_0/IP_IN PAD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm
Xlv_nand_0 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_9178_38525# A lv_nand
Xlv_nand_1 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_1184_38534# PDRV0 lv_nand
X0 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X1 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X2 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_882_55933# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X4 a_882_55933# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X5 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X6 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X7 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X8 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X9 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X10 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X11 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
D0 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D1 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D2 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D3 comp018green_inpath_cms_smt_0/VSUBS w_11000_43887# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D4 A w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
D5 SL w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
X12 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
D6 comp018green_inpath_cms_smt_0/VSUBS PDRV0 diode_pd2nw_03v3 pj=1.92u area=0.2304p
D7 comp018green_inpath_cms_smt_0/VSUBS PDRV1 diode_pd2nw_03v3 pj=1.92u area=0.2304p
X13 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt gf180mcu_ocd_io__bi_a A ANA CS DVDD IE OE PD PDRV0 PDRV1 PU SL VDD Y PAD VSS
+ DVSS
XGF_NI_BI_T_BASE_0 PD IE SL A OE CS PU PDRV0 PDRV1 Y GF_NI_BI_T_BASE_0/ndrive_y_<0>
+ GF_NI_BI_T_BASE_0/ndrive_x_<0> GF_NI_BI_T_BASE_0/ndrive_x_<1> GF_NI_BI_T_BASE_0/ndrive_Y_<1>
+ GF_NI_BI_T_BASE_0/ndrive_x_<2> GF_NI_BI_T_BASE_0/ndrive_y_<2> GF_NI_BI_T_BASE_0/ndrive_x_<3>
+ GF_NI_BI_T_BASE_0/ndrive_Y_<3> GF_NI_BI_T_BASE_0/pdrive_x_<0> GF_NI_BI_T_BASE_0/pdrive_y_<0>
+ GF_NI_BI_T_BASE_0/pdrive_y_<1> GF_NI_BI_T_BASE_0/pdrive_x_<1> GF_NI_BI_T_BASE_0/pdrive_x_<2>
+ GF_NI_BI_T_BASE_0/pdrive_y_<2> GF_NI_BI_T_BASE_0/pdrive_y_<3> GF_NI_BI_T_BASE_0/pdrive_x_<3>
+ VDD VDD DVDD DVDD VDD VDD DVSS VSS DVSS DVSS DVDD DVDD DVDD VSS PAD a_3151_58293#
+ DVDD DVDD DVDD DVDD DVDD DVDD VSS ANA DVSS DVSS DVDD DVDD DVDD VDD VSS VDD DVSS
+ DVDD VDD DVSS GF_NI_BI_T_BASE
.ends

.subckt GF_NI_FILL10_1short VSS VDD DVSS DVDD
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0short DVSS DVDD VDD VSS
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1short
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__tiel_4 VDD VNW VPW VSS ZERO
X0 ZERO a_112_319# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_112_319# a_112_319# VDD VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.6072p ps=3.64u w=1.38u l=0.28u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__tieh_4 VDD VNW VPW VSS ONE
X0 a_112_319# a_112_319# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 ONE a_112_319# VDD VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.6072p ps=3.64u w=1.38u l=0.28u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__buff_12 VDD VNW VPW VSS A Y
X0 VSS a_172_68# Y VPW nfet_03v3 ad=0.985p pd=3.97u as=0.26p ps=1.52u w=1u l=0.28u
X1 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 VDD A a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X4 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X5 VDD a_172_68# Y VNW pfet_03v3 ad=1.3593p pd=4.73u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 a_172_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X7 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X9 Y a_172_68# VDD VNW pfet_03v3 ad=0.36915p pd=1.915u as=0.3588p ps=1.9u w=1.38u l=0.28u
X10 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X11 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X14 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X16 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X18 VSS A a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X19 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X20 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.2675p ps=1.535u w=1u l=0.28u
X21 VDD A a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X22 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X24 a_172_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X25 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X26 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X27 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X28 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X29 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.36915p ps=1.915u w=1.38u l=0.28u
X30 VSS A a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X31 Y a_172_68# VSS VPW nfet_03v3 ad=0.2675p pd=1.535u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt constant_block zero one vdd vss
Xgf180mcu_as_sc_mcu7t3v3__fillcap_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__fillcap_4
Xgf180mcu_as_sc_mcu7t3v3__fillcap_4_1 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__fillcap_4
Xgf180mcu_as_sc_mcu7t3v3__tiel_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_0/A
+ gf180mcu_as_sc_mcu7t3v3__tiel_4
Xgf180mcu_as_sc_mcu7t3v3__tieh_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_1/A
+ gf180mcu_as_sc_mcu7t3v3__tieh_4
Xgf180mcu_as_sc_mcu7t3v3__buff_12_1 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_1/A
+ one gf180mcu_as_sc_mcu7t3v3__buff_12
Xgf180mcu_as_sc_mcu7t3v3__buff_12_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_0/A
+ zero gf180mcu_as_sc_mcu7t3v3__buff_12
.ends

.subckt gf180mcu_ocd_io__fill10x VDD one zero DVDD DVSS VSS
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0short
Xconstant_block_0 zero one VDD VSS constant_block
.ends

.subckt comp018green_esd_rc_v5p0 VRC VPLUS VMINUS
X0 a_353_2269# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X1 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_353_3389# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X3 a_353_2829# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X4 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_353_1709# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X6 a_353_1709# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X7 a_353_2829# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X8 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X9 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X10 VRC a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X11 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X12 a_353_1149# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X13 VPLUS a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X14 a_353_2269# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X15 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X16 a_353_3389# a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X17 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X18 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X19 a_353_1149# a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
.ends

.subckt nmos_clamp_20_50_4_DVSS a_582_632# w_n51_n51# a_1237_1481#
X0 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_DVSS comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VMINUS
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0
Xnmos_clamp_20_50_4_DVSS_0 comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
+ a_4685_27917# nmos_clamp_20_50_4_DVSS
X0 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X10 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X11 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X25 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X33 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X39 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt GF_NI_DVSS_BASE DVDD m2_2292_38400# a_12742_47643# DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
Xcomp018green_esd_clamp_v5p0_DVSS_0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ DVSS comp018green_esd_clamp_v5p0_DVSS
D0 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
D1 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D2 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D3 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X1 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
X2 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
X3 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__dvss DVDD DVSS VDD VSS
XGF_NI_DVSS_BASE_0 DVDD VDD VSS DVSS DVDD GF_NI_DVSS_BASE
.ends

.subckt comp018green_esd_hbm w_n51_7356# a_1131_1121# dw_n51_n51#
D0 dw_n51_n51# a_1131_1121# diode_nd2ps_06v0 pj=0.106m area=0.15n
D1 dw_n51_n51# a_1131_1121# diode_nd2ps_06v0 pj=0.106m area=0.15n
D2 a_1131_1121# w_n51_7356# diode_pd2nw_06v0 pj=0.106m area=0.15n
D3 dw_n51_n51# a_1131_1121# diode_nd2ps_06v0 pj=0.106m area=0.15n
D4 dw_n51_n51# a_1131_1121# diode_nd2ps_06v0 pj=0.106m area=0.15n
D5 a_1131_1121# w_n51_7356# diode_pd2nw_06v0 pj=0.106m area=0.15n
D6 a_1131_1121# w_n51_7356# diode_pd2nw_06v0 pj=0.106m area=0.15n
D7 a_1131_1121# w_n51_7356# diode_pd2nw_06v0 pj=0.106m area=0.15n
.ends

.subckt GF_NI_ASIG_5P0_BASE a_13985_889# m2_828_38097# comp018green_esd_hbm_0/a_1131_1121#
+ m2_13160_36497# w_1350_806# w_2400_15668#
Xcomp018green_esd_hbm_0 w_2400_15668# comp018green_esd_hbm_0/a_1131_1121# w_1350_806#
+ comp018green_esd_hbm
X0 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X1 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X2 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X3 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X4 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X5 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X6 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X7 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X8 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X9 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X10 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X11 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X12 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X13 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X14 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X15 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X16 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X17 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X18 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X19 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X20 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X21 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X22 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X23 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X24 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X25 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X26 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X27 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X28 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X29 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
D0 w_1350_806# w_2400_15668# diode_nd2ps_06v0 pj=82u area=40p
X30 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X31 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X32 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
D1 w_1350_806# w_2400_15668# diode_nd2ps_06v0 pj=82u area=40p
X33 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
D2 w_1350_806# w_2400_15668# diode_nd2ps_06v0 pj=82u area=40p
X34 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
X35 w_2400_15668# w_1350_806# cap_nmos_06v0 c_width=15u c_length=15u
D3 w_1350_806# w_2400_15668# diode_nd2ps_06v0 pj=82u area=40p
.ends

.subckt gf180mcu_ocd_io__asig_5p0 DVDD DVSS VDD ASIG5V VSS
XGF_NI_ASIG_5P0_BASE_0 VSS VDD ASIG5V VSS DVSS DVDD GF_NI_ASIG_5P0_BASE
.ends

.subckt nmos_clamp_20_50_4_DVDD a_582_632# w_n51_n51# a_1237_1481#
X0 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_DVDD comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VMINUS
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0
Xnmos_clamp_20_50_4_DVDD_0 comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
+ a_4685_27917# nmos_clamp_20_50_4_DVDD
X0 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X10 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X11 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X25 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X33 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X39 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt GF_NI_DVDD_BASE DVSS a_246_47643# a_13001_27179# m2_2279_36800# comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS
+ DVDD
Xcomp018green_esd_clamp_v5p0_DVDD_0 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS
+ comp018green_esd_clamp_v5p0_DVDD
D0 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
X0 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
D1 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
D2 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
D3 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
X1 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
X2 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
X3 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__dvdd DVSS VDD VSS DVDD
XGF_NI_DVDD_BASE_0 DVSS VSS VSS VSS DVSS DVDD GF_NI_DVDD_BASE
.ends

.subckt GF_NI_IN_S_BASE PD PU Y ndrive_y_<0> ndrive_x_<0> ndrive_x_<1> ndrive_Y_<1>
+ ndrive_x_<2> ndrive_y_<2> ndrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_y_<0> pdrive_y_<1>
+ pdrive_x_<1> pdrive_x_<2> pdrive_y_<2> pdrive_y_<3> pdrive_x_<3> m3_1771_39126#
+ w_11000_43887# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ m2_1886_52816# comp018green_inpath_cms_smt_0/m3_9619_4882# w_835_53274# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_esd_cdm_0/w_454_3720# m3_10025_37504# PAD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ a_12390_41548# m1_3608_46684# comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ tie_poly_res_0/VSUBS comp018green_sigbuf_1_0/DVSS comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_sigbuf_1_0/DVDD comp018green_inpath_cms_smt_0/m1_10570_5335# comp018green_inpath_cms_smt_0/VSUBS
+ w_11042_41027# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_predrv_3/DVDD w_13720_39292# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
Xlv_nand_2 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_5236_36986# w_13720_39292#
+ lv_nand
Xlv_nand_3 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_4812_38523# w_11184_44921#
+ lv_nand
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ pdrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> comp018green_out_predrv_3/DVDD
+ ndrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ ndrive_y_<2> pdrive_y_<2> pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ ndrive_y_<0> pdrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ ndrive_x_<2> pdrive_x_<1> PAD ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_out_paddrv_16T
Xtie_poly_res_0 w_11184_44921# comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS
+ w_835_53274# tie_poly_res
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/DVSS comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/ZB m1_9774_36986# m1_9537_37107# comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<0> pdrive_y_<0> pdrive_x_<0> comp018green_out_predrv_0/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD m1_9174_38525# m1_9257_38818# comp018green_out_sigbuf_a
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<2> pdrive_y_<2> pdrive_x_<2> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<3> pdrive_y_<3> pdrive_x_<3> comp018green_out_predrv_1/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_0/EN m1_1178_38534# m1_1183_38806#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<1> pdrive_y_<1> pdrive_x_<1> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/CS
+ PU comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/CS
+ w_11000_43887# m1_3608_46684# comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/m3_9619_4882#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
+ Y comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/m1_10570_5335#
+ comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484# PD w_835_53274#
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_1/EN m1_5236_36986# m1_5084_37107#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_sigbuf_oe_1 comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/EN m1_4812_38523# m1_4626_36747#
+ comp018green_out_sigbuf_oe
Xlv_inv_0 w_13720_39292# m1_1183_38806# m1_1178_38534# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_1 w_13720_39292# m1_9257_38818# m1_9174_38525# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_2 w_13720_39292# m1_9537_37107# m1_9774_36986# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_3 w_13720_39292# m1_4626_36747# m1_4812_38523# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_4 w_13720_39292# m1_9774_36986# w_11184_44921# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_6 w_13720_39292# m1_5084_37107# m1_5236_36986# tie_poly_res_0/VSUBS lv_inv
Xcomp018green_esd_cdm_0 comp018green_esd_cdm_0/IP_IN PAD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm
Xlv_nand_0 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_9174_38525# w_11184_44921#
+ lv_nand
Xlv_nand_1 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_1178_38534# w_11184_44921#
+ lv_nand
X0 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X1 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X2 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X4 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X5 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X6 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X7 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X8 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X9 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
D0 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D1 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D2 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D3 comp018green_inpath_cms_smt_0/VSUBS w_11000_43887# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D4 w_11184_44921# w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
D5 w_11184_44921# w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
X10 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
D6 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D7 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
X11 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt gf180mcu_ocd_io__in_s DVDD PD PU VDD Y PAD VSS DVSS
XGF_NI_IN_S_BASE_0 PD PU Y GF_NI_IN_S_BASE_0/ndrive_y_<0> GF_NI_IN_S_BASE_0/ndrive_x_<0>
+ GF_NI_IN_S_BASE_0/ndrive_x_<1> GF_NI_IN_S_BASE_0/ndrive_Y_<1> GF_NI_IN_S_BASE_0/ndrive_x_<2>
+ GF_NI_IN_S_BASE_0/ndrive_y_<2> GF_NI_IN_S_BASE_0/ndrive_x_<3> GF_NI_IN_S_BASE_0/ndrive_Y_<3>
+ GF_NI_IN_S_BASE_0/pdrive_x_<0> GF_NI_IN_S_BASE_0/pdrive_y_<0> GF_NI_IN_S_BASE_0/pdrive_y_<1>
+ GF_NI_IN_S_BASE_0/pdrive_x_<1> GF_NI_IN_S_BASE_0/pdrive_x_<2> GF_NI_IN_S_BASE_0/pdrive_y_<2>
+ GF_NI_IN_S_BASE_0/pdrive_y_<3> GF_NI_IN_S_BASE_0/pdrive_x_<3> VDD VDD DVDD DVDD
+ DVSS VDD VDD DVSS VSS DVSS DVSS DVDD DVDD DVDD VSS PAD DVDD DVDD DVDD DVDD DVDD
+ DVDD VSS DVSS DVSS DVDD DVDD VDD VSS VDD DVSS DVDD VDD DVSS GF_NI_IN_S_BASE
.ends

.subckt GF_NI_VSS_BASE DVSS DVDD VDD m3_12861_12842# m3_7265_24036# m3_7265_54442#
+ m3_5168_44842# m3_9927_40042# m3_12297_28842# m3_7874_12842# m3_4851_11242# m3_7265_20836#
+ m3_7265_43242# m3_12297_24036# m3_12297_54442# m3_7265_41642# m3_4851_17636# m3_10244_48042#
+ m3_12297_20836# m3_2481_11242# m3_12297_43242# m3_12861_33636# m3_9927_28842# m3_12861_1636#
+ m3_12297_41642# m3_10244_44842# m3_2481_17636# m3_5168_1636# m3_12861_56043# m3_2798_27242#
+ m3_7874_33636# m3_9927_24036# m3_9927_54442# m3_7874_56043# m3_4851_30436# m3_7874_1636#
+ m3_9927_20836# m3_9927_43242# m3_2798_1636# m3_9927_41642# m3_7265_46442# m3_2798_12842#
+ m3_2481_30436# m3_7265_14436# m3_4851_40042# m3_5168_27242# m3_12861_8036# m3_5168_8036#
+ m3_12297_46442# m3_12861_4836# m3_12297_14436# m3_5168_4836# m3_2481_40042# m3_7874_8036#
+ m2_2292_38400# m3_12861_48042# m3_2798_8036# m3_4851_28842# m3_2798_33636# m3_5168_12842#
+ m3_7874_4836# m3_10244_1636# m3_9927_46442# m3_12861_44842# m3_7874_48042# m3_2798_56043#
+ m3_10244_27242# m3_4851_24036# m3_7265_11242# m3_2798_4836# m3_4851_54442# m3_9927_14436#
+ m3_2481_28842# m3_7874_44842# m3_7265_17636# m3_4851_20836# m3_4851_43242# m3_12297_11242#
+ m3_2481_24036# m3_2481_54442# m3_4851_41642# m3_5168_33636# m3_10244_12842# m3_12297_17636#
+ m3_2481_20836# m3_2481_43242# m3_10244_8036# m3_5168_56043# m3_2481_41642# m3_7265_30436#
+ m3_9927_11242# m3_10244_4836# m3_9927_17636# m3_2798_48042# m3_12297_30436# m3_10244_33636#
+ m3_7265_40042# m3_4851_46442# m3_2798_44842# m3_12861_27242# m3_10244_56043# m3_4851_14436#
+ VSS m3_12297_40042# m3_7874_27242# m3_2481_46442# comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ m3_9927_30436# m3_2481_14436# m3_7265_28842# m3_5168_48042#
Xcomp018green_esd_clamp_v5p0_DVSS_0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ VSS comp018green_esd_clamp_v5p0_DVSS
D0 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
D1 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D2 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D3 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X1 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
X2 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
X3 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__vss DVDD VDD VSS DVSS
XGF_NI_VSS_BASE_0 DVSS DVDD VDD DVSS DVDD DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVDD
+ DVDD DVDD DVDD DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVSS DVDD DVSS DVDD DVSS DVSS
+ DVSS DVSS DVDD DVDD DVSS DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVDD
+ DVSS DVSS DVSS DVDD DVSS DVDD DVSS DVDD DVSS VDD DVSS DVSS DVDD DVSS DVSS DVSS DVSS
+ DVDD DVSS DVSS DVSS DVSS DVDD DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVDD DVDD DVDD
+ DVDD DVDD DVDD DVSS DVSS DVDD DVDD DVDD DVSS DVSS DVDD DVDD DVDD DVSS DVDD DVSS
+ DVDD DVSS DVDD DVDD DVSS DVSS DVSS DVDD VSS DVDD DVSS DVDD VDD DVDD DVDD DVDD DVSS
+ GF_NI_VSS_BASE
.ends

.subckt moscap_corner_1 a_5519_6541# a_5519_529# a_4904_32#
X0 a_5519_529# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X1 a_5519_6541# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X2 a_5519_529# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X3 a_5519_6541# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt moscap_corner VMINUS a_647_6541# a_647_529#
X0 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X6 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X7 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt nmos_clamp_20_50_4 a_582_632# w_n51_n51# a_1237_1481#
X0 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_rc_v5p0_1 VRC VPLUS VMINUS
X0 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_n2894_17198# a_n2614_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X5 a_n1774_17198# a_n2054_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X6 a_n1214_17198# a_n1494_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X7 a_n2894_17198# a_n3174_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X8 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X9 a_n2334_17198# a_n2614_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X10 a_n1214_17198# a_n934_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X11 a_n3454_17198# VPLUS VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X12 a_n1774_17198# a_n1494_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X13 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X14 a_n2334_17198# a_n2054_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X15 a_n654_17198# a_n934_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X16 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X17 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X18 a_n3454_17198# a_n3174_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X19 a_n654_17198# VRC VPLUS ppolyf_u r_width=0.8u r_length=63.855u
.ends

.subckt comp018green_esd_clamp_v5p0_1 top_route_0/VSUBS comp018green_esd_rc_v5p0_1_0/VPLUS
Xnmos_clamp_20_50_4_0 top_route_0/VSUBS comp018green_esd_rc_v5p0_1_0/VPLUS a_4685_27789#
+ nmos_clamp_20_50_4
Xcomp018green_esd_rc_v5p0_1_0 comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS
+ top_route_0/VSUBS comp018green_esd_rc_v5p0_1
X0 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 comp018green_esd_rc_v5p0_1_0/VPLUS a_2805_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X11 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X25 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X38 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X39 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_2 comp018green_esd_rc_v5p0_0/VPLUS top_route_1_0/VSUBS
Xnmos_clamp_20_50_4_0 top_route_1_0/VSUBS comp018green_esd_rc_v5p0_0/VPLUS a_4685_27789#
+ nmos_clamp_20_50_4
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ top_route_1_0/VSUBS comp018green_esd_rc_v5p0
X0 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X11 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X25 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X38 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X39 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt ESD_CLAMP_COR power_via_cor_3_0/m1_14757_49610# power_via_cor_5_0/m1_14757_35210#
+ power_via_cor_5_0/m1_14757_49610# comp018green_esd_clamp_v5p0_1_0/comp018green_esd_rc_v5p0_1_0/VPLUS
+ power_via_cor_3_0/m1_14757_35210# VSUBS comp018green_esd_clamp_v5p0_2_0/comp018green_esd_rc_v5p0_0/VPLUS
Xcomp018green_esd_clamp_v5p0_1_0 VSUBS comp018green_esd_clamp_v5p0_1_0/comp018green_esd_rc_v5p0_1_0/VPLUS
+ comp018green_esd_clamp_v5p0_1
Xcomp018green_esd_clamp_v5p0_2_0 comp018green_esd_clamp_v5p0_2_0/comp018green_esd_rc_v5p0_0/VPLUS
+ VSUBS comp018green_esd_clamp_v5p0_2
.ends

.subckt moscap_corner_2 VMINUS a_647_6541# a_5519_529#
X0 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_5519_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_5519_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt moscap_corner_3 VMINUS a_7955_529# a_3083_6541#
X0 a_7955_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt GF_NI_COR_BASE ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_35210# ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_49610#
+ ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_35210# moscap_corner_0/a_647_6541# moscap_corner_6/a_647_529#
+ VDD ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_49610# moscap_corner_6/a_647_6541#
+ moscap_corner_4/a_647_529# moscap_corner_0/a_647_529# DVDD VSS moscap_corner_4/a_647_6541#
+ moscap_corner_1/a_647_529#
Xmoscap_corner_1_0 moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# VSS moscap_corner_1
Xmoscap_corner_0 VSS moscap_corner_0/a_647_6541# moscap_corner_0/a_647_529# moscap_corner
Xmoscap_corner_1 VSS moscap_corner_1/a_647_529# moscap_corner_1/a_647_529# moscap_corner
Xmoscap_corner_2 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner
Xmoscap_corner_3 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
Xmoscap_corner_5 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
Xmoscap_corner_4 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner
Xmoscap_corner_6 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
XESD_CLAMP_COR_0 ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_49610# ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_35210#
+ ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_49610# VDD ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_35210#
+ VSS DVDD ESD_CLAMP_COR
Xmoscap_corner_2_0 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner_2
Xmoscap_corner_3_0 VSS moscap_corner_1/a_647_529# moscap_corner_1/a_647_529# moscap_corner_3
.ends

.subckt gf180mcu_ocd_io__cor VDD DVDD VSS
XGF_NI_COR_BASE_0 VSS VSS VSS DVDD DVDD VDD VSS DVDD DVDD DVDD DVDD VSS DVDD DVDD
+ GF_NI_COR_BASE
.ends

.subckt GF_NI_VDD_BASE DVSS DVDD VSS m3_9927_12842# m3_7265_56043# m3_5168_14436#
+ m3_7265_52842# m3_12297_33636# m3_2798_11242# m3_12297_56043# m3_2798_17636# m3_9927_1636#
+ m3_12297_52842# m3_7265_8036# m3_12861_28842# m3_9927_33636# m3_7265_4836# m3_7874_28842#
+ m3_12861_24036# m3_12861_54442# m3_10244_14436# m3_4851_27242# m3_9927_56043# m3_5168_11242#
+ m3_9927_52842# m3_7874_24036# m3_7874_54442# m3_2798_30436# m3_12861_20836# m3_12861_43242#
+ m3_5168_17636# m3_12861_41642# m3_7265_48042# m3_2481_27242# m3_7874_20836# m3_9927_8036#
+ m3_7874_43242# m3_12297_1636# m3_7874_41642# m3_4851_12842# m3_7265_44842# m3_9927_4836#
+ m3_12297_48042# m3_10244_11242# m3_5168_30436# m3_2481_12842# m3_12297_44842# m3_10244_17636#
+ m3_2481_1636# m3_2798_28842# m3_9927_48042# m3_4851_33636# m3_12297_8036# m3_12861_14436#
+ m3_2798_24036# m3_2798_54442# m3_4851_56043# m3_9927_44842# m3_12297_4836# m3_4851_52842#
+ m3_7874_14436# m3_2481_33636# m3_10244_30436# m3_2798_20836# m3_2798_43242# m3_2798_41642#
+ m3_4851_1636# m3_2481_56043# m3_5168_28842# m3_2481_8036# m3_2481_52842# m3_7265_27242#
+ m3_5168_24036# m3_2481_4836# m3_5168_54442# m3_12861_11242# m3_5168_20836# m3_5168_43242#
+ m3_12297_27242# m3_12861_17636# m3_7874_11242# m3_5168_41642# m3_4851_8036# m3_10244_28842#
+ m3_4851_48042# m3_7265_12842# m3_7874_17636# m3_4851_4836# m3_10244_24036# m3_2798_14436#
+ m3_10244_54442# m3_4851_44842# m3_9927_27242# m3_12297_12842# m3_2481_48042# VDD
+ m3_12861_30436# m3_10244_20836# m3_10244_43242# m3_7265_1636# m3_10244_41642# m3_2481_44842#
+ m3_7874_30436# m3_7265_33636#
Xcomp018green_esd_clamp_v5p0_DVDD_0 VDD VSS comp018green_esd_clamp_v5p0_DVDD
D0 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X0 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
D1 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D2 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D3 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X1 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
X2 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
X3 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__vdd DVDD DVSS VDD VSS
XGF_NI_VDD_BASE_0 DVSS DVDD VSS DVSS DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVSS
+ DVSS DVDD DVSS DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVDD
+ DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVSS DVDD DVDD
+ DVSS DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVDD DVDD DVDD DVSS DVSS DVSS DVSS DVDD
+ DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVSS DVSS DVDD DVSS DVDD DVDD DVDD
+ DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVSS DVSS
+ DVSS DVSS VDD DVDD DVDD DVDD DVSS DVDD DVSS DVDD DVSS GF_NI_VDD_BASE
.ends

.subckt chip_half_frame DVDD analog_PAD[0] analog_PAD[1] analog_PAD[2] analog_PAD[3]
+ input_PAD[0] input_PAD[1] input_PAD[2] input_PAD[3] clk_PAD rst_n_PAD bidir_PAD[0]
+ bidir_PAD[1] bidir_PAD[2] bidir_PAD[3] bidir_PAD[4] bidir_PAD[5] bidir_PAD[6] bidir_PAD[7]
+ bidir_PAD[8] bidir_PAD[9] bidir_PAD[10] bidir_PAD[11] bidir_PAD[12] bidir_PAD[13]
+ bidir_PAD[14] bidir_PAD[15] bidir_PAD[16] bidir_PAD[17] bidir_PAD[18] bidir_PAD[19]
+ bidir_PAD[20] bidir_PAD[21] bidir_PAD[22] bidir_PAD[23] bidir_PAD[24] bidir_PAD[25]
+ bidir_PAD[26] bidir_PAD[27] bidir_PAD[28] bidir_PAD[29] bidir_PAD[30] bidir_PAD[31]
+ bidir_PAD[32] bidir_PAD[33] bidir_PAD[34] bidir_PAD[35] bidir_PAD[36] bidir_PAD[37]
+ bidir_PAD[38] bidir_PAD[39] bidir_PAD[40] bidir_PAD[41] bidir_PAD[42] bidir_PAD[43]
+ bidir_PAD[44] bidir_PAD[45] gf180mcu_ocd_io__fill10x_47/one gf180mcu_ocd_io__bi_a_15/SL
+ gf180mcu_ocd_io__bi_a_38/PD gf180mcu_ocd_io__bi_a_16/IE gf180mcu_ocd_io__bi_a_43/PD
+ gf180mcu_ocd_io__bi_a_0/PD gf180mcu_ocd_io__bi_a_8/IE gf180mcu_ocd_io__bi_a_16/PD
+ gf180mcu_ocd_io__fill10x_59/zero gf180mcu_ocd_io__bi_a_18/PDRV0 gf180mcu_ocd_io__bi_a_35/PD
+ gf180mcu_ocd_io__bi_a_19/IE gf180mcu_ocd_io__bi_a_11/Y gf180mcu_ocd_io__bi_a_1/Y
+ gf180mcu_ocd_io__bi_a_40/PD gf180mcu_ocd_io__bi_a_8/PD gf180mcu_ocd_io__bi_a_17/A
+ gf180mcu_ocd_io__bi_a_13/OE gf180mcu_ocd_io__bi_a_27/PD gf180mcu_ocd_io__bi_a_19/PD
+ gf180mcu_ocd_io__fill10x_271/one gf180mcu_ocd_io__bi_a_32/PD gf180mcu_ocd_io__bi_a_15/PDRV0
+ gf180mcu_ocd_io__bi_a_4/OE gf180mcu_ocd_io__bi_a_15/OE gf180mcu_ocd_io__bi_a_10/OE
+ gf180mcu_ocd_io__bi_a_24/PD gf180mcu_ocd_io__fill10x_287/zero gf180mcu_ocd_io__bi_a_16/PDRV0
+ gf180mcu_ocd_io__fill10x_350/one gf180mcu_ocd_io__bi_a_42/Y gf180mcu_ocd_io__bi_a_17/Y
+ gf180mcu_ocd_io__fill10x_323/one gf180mcu_ocd_io__bi_a_13/PD gf180mcu_ocd_io__bi_a_5/PDRV0
+ gf180mcu_ocd_io__bi_a_5/PDRV1 gf180mcu_ocd_io__in_c_2/Y gf180mcu_ocd_io__fill10x_65/zero
+ gf180mcu_ocd_io__fill10x_395/one gf180mcu_ocd_io__bi_a_7/PDRV1 gf180mcu_ocd_io__bi_a_33/A
+ gf180mcu_ocd_io__fill10x_190/one gf180mcu_ocd_io__fill10x_264/zero gf180mcu_ocd_io__fill10x_94/one
+ gf180mcu_ocd_io__bi_a_7/SL gf180mcu_ocd_io__bi_a_10/PD gf180mcu_ocd_io__bi_a_45/IE
+ gf180mcu_ocd_io__bi_a_14/PDRV1 gf180mcu_ocd_io__bi_a_9/PDRV0 gf180mcu_ocd_io__bi_a_9/SL
+ gf180mcu_ocd_io__bi_a_13/Y gf180mcu_ocd_io__bi_a_37/IE gf180mcu_ocd_io__fill10x_47/zero
+ gf180mcu_ocd_io__bi_a_42/IE gf180mcu_ocd_io__bi_a_6/A gf180mcu_ocd_io__bi_a_40/PDRV1
+ gf180mcu_ocd_io__bi_a_43/Y gf180mcu_ocd_io__bi_a_29/IE gf180mcu_ocd_io__bi_a_36/A
+ gf180mcu_ocd_io__fill10_310x/zero gf180mcu_ocd_io__bi_a_16/A gf180mcu_ocd_io__bi_a_34/IE
+ gf180mcu_ocd_io__bi_a_10/A gf180mcu_ocd_io__bi_a_7/OE gf180mcu_ocd_io__bi_a_26/IE
+ gf180mcu_ocd_io__bi_a_21/SL gf180mcu_ocd_io__fill10x_258/one gf180mcu_ocd_io__bi_a_9/OE
+ gf180mcu_ocd_io__bi_a_31/IE gf180mcu_ocd_io__fill10x_341/zero gf180mcu_ocd_io__bi_a_40/PDRV0
+ gf180mcu_ocd_io__fill10x_102/zero gf180mcu_ocd_io__bi_a_41/PDRV1 gf180mcu_ocd_io__bi_a_23/IE
+ gf180mcu_ocd_io__bi_a_4/PDRV0 gf180mcu_ocd_io__bi_a_6/Y gf180mcu_ocd_io__in_s_0/Y
+ gf180mcu_ocd_io__bi_a_16/Y gf180mcu_ocd_io__fill10x_307/one gf180mcu_ocd_io__bi_a_35/A
+ gf180mcu_ocd_io__fill10x_401/one gf180mcu_ocd_io__bi_a_45/SL gf180mcu_ocd_io__bi_a_39/PU
+ gf180mcu_ocd_io__fill10x_126/zero gf180mcu_ocd_io__bi_a_44/PU gf180mcu_ocd_io__bi_a_6/PDRV0
+ gf180mcu_ocd_io__bi_a_41/PDRV0 gf180mcu_ocd_io__fill10x_177/one gf180mcu_ocd_io__in_c_4/Y
+ gf180mcu_ocd_io__bi_a_1/IE gf180mcu_ocd_io__bi_a_21/OE gf180mcu_ocd_io__bi_a_37/SL
+ gf180mcu_ocd_io__bi_a_42/PDRV1 gf180mcu_ocd_io__bi_a_12/IE gf180mcu_ocd_io__fill10x_280/zero
+ gf180mcu_ocd_io__bi_a_42/SL gf180mcu_ocd_io__bi_a_15/IE gf180mcu_ocd_io__fill10x_58/one
+ gf180mcu_ocd_io__bi_a_36/PU gf180mcu_ocd_io__bi_a_1/PD gf180mcu_ocd_io__bi_a_1/SL
+ gf180mcu_ocd_io__bi_a_41/PU gf180mcu_ocd_io__bi_a_42/A gf180mcu_ocd_io__fill10x_36/zero
+ gf180mcu_ocd_io__fill10x_25/one gf180mcu_ocd_io__bi_a_29/SL gf180mcu_ocd_io__bi_a_6/IE
+ gf180mcu_ocd_io__bi_a_8/PDRV0 gf180mcu_ocd_io__bi_a_34/SL gf180mcu_ocd_io__bi_a_15/PD
+ gf180mcu_ocd_io__bi_a_28/PU gf180mcu_ocd_io__bi_a_21/IE gf180mcu_ocd_io__bi_a_38/CS
+ gf180mcu_ocd_io__bi_a_33/PU gf180mcu_ocd_io__bi_a_6/PD gf180mcu_ocd_io__bi_a_43/CS
+ gf180mcu_ocd_io__bi_a_42/PDRV0 gf180mcu_ocd_io__bi_a_12/A gf180mcu_ocd_io__bi_a_26/SL
+ gf180mcu_ocd_io__fill10x_103/one gf180mcu_ocd_io__bi_a_21/PD gf180mcu_ocd_io__bi_a_43/PDRV1
+ gf180mcu_ocd_io__bi_a_3/A gf180mcu_ocd_io__bi_a_31/SL gf180mcu_ocd_io__bi_a_7/PDRV0
+ gf180mcu_ocd_io__bi_a_25/PU gf180mcu_ocd_io__bi_a_38/A gf180mcu_ocd_io__fill10x_54/one
+ gf180mcu_ocd_io__bi_a_35/CS gf180mcu_ocd_io__bi_a_30/PU gf180mcu_ocd_io__bi_a_40/CS
+ gf180mcu_ocd_io__bi_a_23/SL gf180mcu_ocd_io__in_c_3/PU gf180mcu_ocd_io__bi_a_27/CS
+ gf180mcu_ocd_io__bi_a_1/OE gf180mcu_ocd_io__bi_a_22/PU gf180mcu_ocd_io__fill10x_355/zero
+ gf180mcu_ocd_io__bi_a_3/PDRV0 gf180mcu_ocd_io__bi_a_17/SL gf180mcu_ocd_io__bi_a_32/CS
+ gf180mcu_ocd_io__fill10x_163/one gf180mcu_ocd_io__bi_a_43/PDRV0 gf180mcu_ocd_io__in_c_0/Y
+ gf180mcu_ocd_io__bi_a_45/OE gf180mcu_ocd_io__bi_a_44/PDRV1 gf180mcu_ocd_io__bi_a_24/CS
+ gf180mcu_ocd_io__fill10x_287/one gf180mcu_ocd_io__bi_a_0/PDRV1 gf180mcu_ocd_io__bi_a_2/PDRV0
+ gf180mcu_ocd_io__bi_a_3/Y gf180mcu_ocd_io__bi_a_37/OE gf180mcu_ocd_io__bi_a_12/SL
+ gf180mcu_ocd_io__bi_a_19/A gf180mcu_ocd_io__bi_a_42/OE gf180mcu_ocd_io__bi_a_31/A
+ gf180mcu_ocd_io__bi_a_16/PDRV1 gf180mcu_ocd_io__bi_a_11/PU gf180mcu_ocd_io__fill10x_113/zero
+ gf180mcu_ocd_io__bi_a_29/OE gf180mcu_ocd_io__bi_a_8/PDRV1 gf180mcu_ocd_io__bi_a_44/PDRV0
+ gf180mcu_ocd_io__bi_a_44/A gf180mcu_ocd_io__bi_a_34/OE gf180mcu_ocd_io__bi_a_1/PDRV0
+ gf180mcu_ocd_io__fill10x_345/one gf180mcu_ocd_io__bi_a_17/OE gf180mcu_ocd_io__bi_a_13/CS
+ gf180mcu_ocd_io__bi_a_19/PDRV1 gf180mcu_ocd_io__bi_a_45/PDRV1 gf180mcu_ocd_io__bi_a_30/PDRV1
+ gf180mcu_ocd_io__fill10x_22/zero gf180mcu_ocd_io__bi_a_26/OE gf180mcu_ocd_io__bi_a_31/OE
+ gf180mcu_ocd_io__bi_a_45/PD gf180mcu_ocd_io__bi_a_10/CS gf180mcu_ocd_io__bi_a_0/PDRV0
+ gf180mcu_ocd_io__fill10x_389/one gf180mcu_ocd_io__bi_a_19/Y gf180mcu_ocd_io__bi_a_23/OE
+ gf180mcu_ocd_io__bi_a_30/PDRV0 gf180mcu_ocd_io__bi_a_45/PDRV0 gf180mcu_ocd_io__bi_a_37/PD
+ gf180mcu_ocd_io__fill10x_318/one gf180mcu_ocd_io__bi_a_42/PD gf180mcu_ocd_io__bi_a_31/PDRV1
+ gf180mcu_ocd_io__bi_a_0/A gf180mcu_ocd_io__bi_a_28/A gf180mcu_ocd_io__in_c_3/PD
+ gf180mcu_ocd_io__bi_a_29/PD gf180mcu_ocd_io__bi_a_34/PD gf180mcu_ocd_io__fill10x_395/zero
+ gf180mcu_ocd_io__bi_a_6/SL gf180mcu_ocd_io__bi_a_12/OE gf180mcu_ocd_io__bi_a_16/SL
+ gf180mcu_ocd_io__bi_a_26/PD gf180mcu_ocd_io__fill10x_78/one gf180mcu_ocd_io__bi_a_31/PDRV0
+ gf180mcu_ocd_io__fill10x_331/zero gf180mcu_ocd_io__bi_a_31/PD gf180mcu_ocd_io__bi_a_32/PDRV1
+ gf180mcu_ocd_io__bi_a_23/PD gf180mcu_ocd_io__bi_a_0/Y gf180mcu_ocd_io__bi_a_18/A
+ gf180mcu_ocd_io__fill10x_264/one gf180mcu_ocd_io__fill10x_163/zero gf180mcu_ocd_io__fill10x_247/zero
+ gf180mcu_ocd_io__bi_a_2/IE gf180mcu_ocd_io__fill10x_205/zero gf180mcu_ocd_io__fill10x_0/zero
+ gf180mcu_ocd_io__bi_a_32/PDRV0 gf180mcu_ocd_io__bi_a_6/OE gf180mcu_ocd_io__bi_a_18/IE
+ gf180mcu_ocd_io__bi_a_2/PD gf180mcu_ocd_io__bi_a_33/PDRV1 gf180mcu_ocd_io__bi_a_16/OE
+ gf180mcu_ocd_io__fill10x_54/zero gf180mcu_ocd_io__bi_a_4/IE gf180mcu_ocd_io__bi_a_18/PD
+ gf180mcu_ocd_io__bi_a_12/PD gf180mcu_ocd_io__fill10x_294/one gf180mcu_ocd_io__bi_a_20/IE
+ gf180mcu_ocd_io__bi_a_33/Y gf180mcu_ocd_io__bi_a_4/PD gf180mcu_ocd_io__bi_a_23/A
+ gf180mcu_ocd_io__bi_a_39/IE gf180mcu_ocd_io__bi_a_20/PD gf180mcu_ocd_io__bi_a_45/Y
+ gf180mcu_ocd_io__bi_a_18/Y gf180mcu_ocd_io__bi_a_33/PDRV0 gf180mcu_ocd_io__bi_a_44/IE
+ gf180mcu_ocd_io__fill10x_65/one gf180mcu_ocd_io__bi_a_34/PDRV1 gf180mcu_ocd_io__fill10x_336/zero
+ gf180mcu_ocd_io__in_c_1/Y gf180mcu_ocd_io__fill10x_13/one gf180mcu_ocd_io__bi_a_36/IE
+ gf180mcu_ocd_io__in_c_1/PU gf180mcu_ocd_io__bi_a_41/IE gf180mcu_ocd_io__bi_a_20/PU
+ gf180mcu_ocd_io__bi_a_30/A gf180mcu_ocd_io__in_c_0/PU gf180mcu_ocd_io__bi_a_28/IE
+ gf180mcu_ocd_io__bi_a_3/SL gf180mcu_ocd_io__bi_a_33/IE gf180mcu_ocd_io__bi_a_10/Y
+ gf180mcu_ocd_io__fill10x_121/one gf180mcu_ocd_io__bi_a_34/PDRV0 gf180mcu_ocd_io__bi_a_1/PDRV1
+ gf180mcu_ocd_io__bi_a_21/PU gf180mcu_ocd_io__fill10x_71/one gf180mcu_ocd_io__in_s_0/PU
+ gf180mcu_ocd_io__bi_a_35/PDRV1 gf180mcu_ocd_io__bi_a_25/IE gf180mcu_ocd_io__fill10x_138/zero
+ gf180mcu_ocd_io__bi_a_15/PDRV1 gf180mcu_ocd_io__bi_a_30/IE gf180mcu_ocd_io__bi_a_8/A
+ gf180mcu_ocd_io__fill10x_300/zero gf180mcu_ocd_io__bi_a_37/A gf180mcu_ocd_io__bi_a_6/PDRV1
+ gf180mcu_ocd_io__bi_a_5/A gf180mcu_ocd_io__fill10x_171/one gf180mcu_ocd_io__bi_a_19/PU
+ gf180mcu_ocd_io__bi_a_22/IE gf180mcu_ocd_io__bi_a_20/CS gf180mcu_ocd_io__bi_a_21/PDRV1
+ gf180mcu_ocd_io__fill10x_400/zero gf180mcu_ocd_io__bi_a_35/PDRV0 gf180mcu_ocd_io__bi_a_3/OE
+ gf180mcu_ocd_io__bi_a_35/Y gf180mcu_ocd_io__bi_a_39/SL gf180mcu_ocd_io__bi_a_19/SL
+ gf180mcu_ocd_io__bi_a_36/PDRV1 gf180mcu_ocd_io__bi_a_25/A gf180mcu_ocd_io__bi_a_44/SL
+ gf180mcu_ocd_io__bi_a_38/PU gf180mcu_ocd_io__bi_a_14/PU gf180mcu_ocd_io__bi_a_21/CS
+ gf180mcu_ocd_io__bi_a_43/PU gf180mcu_ocd_io__bi_a_36/SL gf180mcu_ocd_io__bi_a_11/IE
+ gf180mcu_ocd_io__bi_a_8/Y gf180mcu_ocd_io__bi_a_41/SL gf180mcu_ocd_io__bi_a_35/PU
+ gf180mcu_ocd_io__fill10x_341/one gf180mcu_ocd_io__bi_a_20/A gf180mcu_ocd_io__bi_a_45/CS
+ gf180mcu_ocd_io__bi_a_36/PDRV0 gf180mcu_ocd_io__bi_a_5/Y gf180mcu_ocd_io__bi_a_32/A
+ gf180mcu_ocd_io__bi_a_40/PU gf180mcu_ocd_io__bi_a_17/PU gf180mcu_ocd_io__bi_a_28/SL
+ gf180mcu_ocd_io__bi_a_19/CS gf180mcu_ocd_io__in_c_1/PD gf180mcu_ocd_io__bi_a_37/PDRV1
+ gf180mcu_ocd_io__fill10x_350/zero gf180mcu_ocd_io__bi_a_22/PDRV1 gf180mcu_ocd_io__bi_a_33/SL
+ gf180mcu_ocd_io__bi_a_27/PU gf180mcu_ocd_io__bi_a_37/CS gf180mcu_ocd_io__bi_a_12/Y
+ gf180mcu_ocd_io__bi_a_32/PU gf180mcu_ocd_io__bi_a_42/CS gf180mcu_ocd_io__bi_a_19/OE
+ gf180mcu_ocd_io__bi_a_25/SL gf180mcu_ocd_io__bi_a_18/PU gf180mcu_ocd_io__fill10x_361/one
+ gf180mcu_ocd_io__bi_a_14/CS gf180mcu_ocd_io__bi_a_29/CS gf180mcu_ocd_io__bi_a_30/SL
+ gf180mcu_ocd_io__bi_a_24/PU gf180mcu_ocd_io__bi_a_0/SL gf180mcu_ocd_io__bi_a_34/CS
+ gf180mcu_ocd_io__bi_a_37/PDRV0 gf180mcu_ocd_io__bi_a_22/PDRV0 gf180mcu_ocd_io__fill10_310x/one
+ gf180mcu_ocd_io__bi_a_22/SL gf180mcu_ocd_io__fill10x_103/zero gf180mcu_ocd_io__bi_a_38/PDRV1
+ gf180mcu_ocd_io__bi_a_23/PDRV1 gf180mcu_ocd_io__bi_a_20/Y gf180mcu_ocd_io__bi_a_26/CS
+ gf180mcu_ocd_io__bi_a_9/IE gf180mcu_ocd_io__fill10x_154/zero gf180mcu_ocd_io__bi_a_15/PU
+ gf180mcu_ocd_io__bi_a_17/CS gf180mcu_ocd_io__bi_a_31/CS gf180mcu_ocd_io__fill10x_307/zero
+ gf180mcu_ocd_io__bi_a_3/IE gf180mcu_ocd_io__bi_a_39/OE gf180mcu_ocd_io__bi_a_2/A
+ gf180mcu_ocd_io__bi_a_9/PD gf180mcu_ocd_io__bi_a_44/OE gf180mcu_ocd_io__bi_a_40/A
+ gf180mcu_ocd_io__bi_a_13/PU gf180mcu_ocd_io__bi_a_17/IE gf180mcu_ocd_io__bi_a_23/CS
+ gf180mcu_ocd_io__fill10x_25/zero gf180mcu_ocd_io__fill10x_102/one gf180mcu_ocd_io__bi_a_3/PD
+ gf180mcu_ocd_io__fill10x_323/zero gf180mcu_ocd_io__bi_a_16/PU gf180mcu_ocd_io__bi_a_38/PDRV0
+ gf180mcu_ocd_io__bi_a_18/CS gf180mcu_ocd_io__bi_a_23/PDRV0 gf180mcu_ocd_io__bi_a_36/OE
+ gf180mcu_ocd_io__bi_a_11/SL gf180mcu_ocd_io__bi_a_17/PD gf180mcu_ocd_io__bi_a_0/OE
+ gf180mcu_ocd_io__bi_a_41/OE gf180mcu_ocd_io__bi_a_39/PDRV1 gf180mcu_ocd_io__bi_a_24/PDRV1
+ gf180mcu_ocd_io__bi_a_18/SL gf180mcu_ocd_io__bi_a_10/PU gf180mcu_ocd_io__in_c_0/PD
+ gf180mcu_ocd_io__bi_a_28/OE gf180mcu_ocd_io__fill10x_247/one gf180mcu_ocd_io__bi_a_33/OE
+ gf180mcu_ocd_io__bi_a_5/PU gf180mcu_ocd_io__bi_a_15/CS gf180mcu_ocd_io__fill10x_190/zero
+ gf180mcu_ocd_io__fill10x_94/zero gf180mcu_ocd_io__bi_a_12/CS gf180mcu_ocd_io__bi_a_2/Y
+ gf180mcu_ocd_io__in_s_0/PD gf180mcu_ocd_io__bi_a_25/OE gf180mcu_ocd_io__bi_a_14/A
+ gf180mcu_ocd_io__bi_a_24/PDRV0 gf180mcu_ocd_io__bi_a_39/PDRV0 gf180mcu_ocd_io__bi_a_27/A
+ gf180mcu_ocd_io__bi_a_39/PD gf180mcu_ocd_io__bi_a_30/OE gf180mcu_ocd_io__fill10x_389/zero
+ gf180mcu_ocd_io__in_c_2/PU gf180mcu_ocd_io__bi_a_9/PU gf180mcu_ocd_io__bi_a_44/PD
+ gf180mcu_ocd_io__bi_a_25/PDRV1 gf180mcu_ocd_io__bi_a_10/PDRV1 gf180mcu_ocd_io__bi_a_16/CS
+ gf180mcu_ocd_io__fill10x_280/one gf180mcu_ocd_io__bi_a_22/OE gf180mcu_ocd_io__bi_a_18/OE
+ gf180mcu_ocd_io__bi_a_34/A gf180mcu_ocd_io__bi_a_36/PD gf180mcu_ocd_io__bi_a_41/PD
+ gf180mcu_ocd_io__bi_a_11/A gf180mcu_ocd_io__bi_a_2/PDRV1 gf180mcu_ocd_io__bi_a_5/CS
+ gf180mcu_ocd_io__bi_a_25/PDRV0 gf180mcu_ocd_io__bi_a_28/PD gf180mcu_ocd_io__bi_a_10/PDRV0
+ gf180mcu_ocd_io__fill10x_171/zero gf180mcu_ocd_io__bi_a_33/PD gf180mcu_ocd_io__bi_a_18/PDRV1
+ gf180mcu_ocd_io__fill10x_266/zero gf180mcu_ocd_io__fill10x_36/one gf180mcu_ocd_io__bi_a_26/PDRV1
+ gf180mcu_ocd_io__bi_a_29/A gf180mcu_ocd_io__bi_a_11/PDRV1 gf180mcu_ocd_io__bi_a_14/Y
+ gf180mcu_ocd_io__bi_a_4/PDRV1 gf180mcu_ocd_io__bi_a_11/OE gf180mcu_ocd_io__bi_a_9/CS
+ gf180mcu_ocd_io__bi_a_25/PD gf180mcu_ocd_io__bi_a_20/PDRV1 gf180mcu_ocd_io__bi_a_30/PD
+ gf180mcu_ocd_io__fill10x_71/zero gf180mcu_ocd_io__fill10x_126/one gf180mcu_ocd_io__bi_a_26/PDRV0
+ gf180mcu_ocd_io__fill10x_59/one gf180mcu_ocd_io__bi_a_11/PDRV0 gf180mcu_ocd_io__bi_a_4/PU
+ gf180mcu_ocd_io__bi_a_22/PD gf180mcu_ocd_io__bi_a_8/SL gf180mcu_ocd_io__bi_a_27/PDRV1
+ gf180mcu_ocd_io__bi_a_12/PDRV1 gf180mcu_ocd_io__bi_a_5/SL gf180mcu_ocd_io__fill10x_106/one
+ gf180mcu_ocd_io__bi_a_6/PU gf180mcu_ocd_io__fill10x_271/zero gf180mcu_ocd_io__bi_a_43/A
+ gf180mcu_ocd_io__bi_a_4/A gf180mcu_ocd_io__in_c_2/PD gf180mcu_ocd_io__bi_a_44/Y
+ gf180mcu_ocd_io__bi_a_11/PD gf180mcu_ocd_io__bi_a_41/A gf180mcu_ocd_io__bi_a_27/PDRV0
+ gf180mcu_ocd_io__bi_a_12/PDRV0 gf180mcu_ocd_io__bi_a_15/A gf180mcu_ocd_io__bi_a_28/PDRV1
+ gf180mcu_ocd_io__bi_a_13/PDRV1 gf180mcu_ocd_io__bi_a_8/PU gf180mcu_ocd_io__bi_a_13/A
+ gf180mcu_ocd_io__bi_a_4/CS gf180mcu_ocd_io__bi_a_38/IE gf180mcu_ocd_io__bi_a_8/OE
+ gf180mcu_ocd_io__bi_a_43/IE gf180mcu_ocd_io__bi_a_20/SL gf180mcu_ocd_io__bi_a_5/OE
+ gf180mcu_ocd_io__fill10x_58/zero gf180mcu_ocd_io__fill10x_336/one gf180mcu_ocd_io__bi_a_7/PU
+ gf180mcu_ocd_io__bi_a_35/IE gf180mcu_ocd_io__bi_a_6/CS gf180mcu_ocd_io__bi_a_5/IE
+ gf180mcu_ocd_io__bi_a_28/PDRV0 gf180mcu_ocd_io__bi_a_13/PDRV0 gf180mcu_ocd_io__bi_a_40/IE
+ gf180mcu_ocd_io__fill10x_258/zero gf180mcu_ocd_io__fill10x_177/zero gf180mcu_ocd_io__bi_a_4/Y
+ gf180mcu_ocd_io__bi_a_29/PDRV1 gf180mcu_ocd_io__bi_a_7/IE gf180mcu_ocd_io__bi_a_27/IE
+ gf180mcu_ocd_io__fill10x_401/zero gf180mcu_ocd_io__bi_a_15/Y gf180mcu_ocd_io__bi_a_5/PD
+ gf180mcu_ocd_io__bi_a_32/IE gf180mcu_ocd_io__bi_a_14/IE gf180mcu_ocd_io__bi_a_3/PU
+ gf180mcu_ocd_io__fill10x_355/one gf180mcu_ocd_io__bi_a_7/PD gf180mcu_ocd_io__bi_a_8/CS
+ gf180mcu_ocd_io__bi_a_20/OE gf180mcu_ocd_io__bi_a_14/PD gf180mcu_ocd_io__bi_a_24/IE
+ gf180mcu_ocd_io__fill10x_331/one gf180mcu_ocd_io__bi_a_29/PDRV0 gf180mcu_ocd_io__bi_a_2/PU
+ gf180mcu_ocd_io__bi_a_2/SL gf180mcu_ocd_io__bi_a_7/CS gf180mcu_ocd_io__bi_a_45/A
+ gf180mcu_ocd_io__bi_a_45/PU gf180mcu_ocd_io__fill10x_345/zero gf180mcu_ocd_io__fill10x_0/one
+ gf180mcu_ocd_io__bi_a_38/SL gf180mcu_ocd_io__bi_a_13/IE gf180mcu_ocd_io__bi_a_1/PU
+ gf180mcu_ocd_io__bi_a_43/SL gf180mcu_ocd_io__bi_a_3/CS gf180mcu_ocd_io__bi_a_7/A
+ gf180mcu_ocd_io__bi_a_37/PU gf180mcu_ocd_io__bi_a_39/A gf180mcu_ocd_io__bi_a_42/PU
+ gf180mcu_ocd_io__bi_a_9/A gf180mcu_ocd_io__bi_a_35/SL gf180mcu_ocd_io__fill10x_266/one
+ gf180mcu_ocd_io__bi_a_29/PU gf180mcu_ocd_io__bi_a_9/PDRV1 gf180mcu_ocd_io__bi_a_39/CS
+ gf180mcu_ocd_io__bi_a_40/SL gf180mcu_ocd_io__bi_a_32/Y gf180mcu_ocd_io__bi_a_0/PU
+ gf180mcu_ocd_io__bi_a_34/PU gf180mcu_ocd_io__bi_a_2/OE gf180mcu_ocd_io__bi_a_2/CS
+ gf180mcu_ocd_io__fill10x_197/zero gf180mcu_ocd_io__bi_a_44/CS gf180mcu_ocd_io__fill10x_318/zero
+ gf180mcu_ocd_io__bi_a_14/SL gf180mcu_ocd_io__bi_a_22/A gf180mcu_ocd_io__bi_a_3/PDRV1
+ gf180mcu_ocd_io__fill10x_121/zero gf180mcu_ocd_io__bi_a_27/SL VDD gf180mcu_ocd_io__bi_a_32/SL
+ gf180mcu_ocd_io__bi_a_17/PDRV1 gf180mcu_ocd_io__bi_a_26/PU gf180mcu_ocd_io__bi_a_36/CS
+ gf180mcu_ocd_io__fill10x_294/zero gf180mcu_ocd_io__bi_a_20/PDRV0 gf180mcu_ocd_io__bi_a_31/PU
+ gf180mcu_ocd_io__bi_a_10/IE gf180mcu_ocd_io__bi_a_41/CS gf180mcu_ocd_io__fill10x_300/one
+ gf180mcu_ocd_io__bi_a_1/CS gf180mcu_ocd_io__bi_a_24/SL gf180mcu_ocd_io__fill10x_13/zero
+ gf180mcu_ocd_io__bi_a_7/Y gf180mcu_ocd_io__bi_a_28/CS gf180mcu_ocd_io__bi_a_21/A
+ gf180mcu_ocd_io__fill10x_78/zero gf180mcu_ocd_io__bi_a_23/PU gf180mcu_ocd_io__bi_a_9/Y
+ gf180mcu_ocd_io__bi_a_33/CS gf180mcu_ocd_io__bi_a_21/PDRV0 gf180mcu_ocd_io__bi_a_0/CS
+ gf180mcu_ocd_io__bi_a_25/CS gf180mcu_ocd_io__bi_a_14/OE gf180mcu_ocd_io__bi_a_30/CS
+ gf180mcu_ocd_io__fill10x_400/one gf180mcu_ocd_io__bi_a_38/OE gf180mcu_ocd_io__bi_a_13/SL
+ gf180mcu_ocd_io__bi_a_19/PDRV0 gf180mcu_ocd_io__bi_a_43/OE gf180mcu_ocd_io__bi_a_12/PU
+ gf180mcu_ocd_io__bi_a_22/CS gf180mcu_ocd_io__fill10x_361/zero gf180mcu_ocd_io__bi_a_35/OE
+ gf180mcu_ocd_io__fill10x_138/one gf180mcu_ocd_io__bi_a_10/SL gf180mcu_ocd_io__bi_a_40/OE
+ gf180mcu_ocd_io__fill10x_22/one gf180mcu_ocd_io__bi_a_14/PDRV0 gf180mcu_ocd_io__bi_a_34/Y
+ gf180mcu_ocd_io__bi_a_1/A gf180mcu_ocd_io__bi_a_27/OE gf180mcu_ocd_io__bi_a_24/A
+ gf180mcu_ocd_io__bi_a_26/A gf180mcu_ocd_io__bi_a_32/OE gf180mcu_ocd_io__bi_a_11/CS
+ gf180mcu_ocd_io__fill10x_113/one gf180mcu_ocd_io__bi_a_0/IE gf180mcu_ocd_io__bi_a_4/SL
+ gf180mcu_ocd_io__bi_a_17/PDRV0 gf180mcu_ocd_io__fill10x_106/zero gf180mcu_ocd_io__bi_a_24/OE
+ VSS
Xgf180mcu_ocd_io__fill10_219 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_208 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_2 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__in_c_3 DVDD gf180mcu_ocd_io__in_c_3/PD gf180mcu_ocd_io__in_c_3/PU
+ VDD gf180mcu_ocd_io__in_c_3/Y input_PAD[1] VSS VSS gf180mcu_ocd_io__in_c
Xgf180mcu_ocd_io__fill10_391 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_380 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_19 gf180mcu_ocd_io__bi_a_19/A gf180mcu_ocd_io__bi_a_19/ANA
+ gf180mcu_ocd_io__bi_a_19/CS DVDD gf180mcu_ocd_io__bi_a_19/IE gf180mcu_ocd_io__bi_a_19/OE
+ gf180mcu_ocd_io__bi_a_19/PD gf180mcu_ocd_io__bi_a_19/PDRV0 gf180mcu_ocd_io__bi_a_19/PDRV1
+ gf180mcu_ocd_io__bi_a_19/PU gf180mcu_ocd_io__bi_a_19/SL VDD gf180mcu_ocd_io__bi_a_19/Y
+ bidir_PAD[2] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_209 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_3 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__in_c_4 DVDD gf180mcu_ocd_io__in_c_4/PD gf180mcu_ocd_io__in_c_4/PU
+ VDD gf180mcu_ocd_io__in_c_4/Y input_PAD[0] VSS VSS gf180mcu_ocd_io__in_c
Xgf180mcu_ocd_io__fill10_381 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_392 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_370 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_4 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_393 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_360 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_382 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_371 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_247 VDD gf180mcu_ocd_io__fill10x_247/one gf180mcu_ocd_io__fill10x_247/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_258 VDD gf180mcu_ocd_io__fill10x_258/one gf180mcu_ocd_io__fill10x_258/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_5 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_383 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_394 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_372 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_180 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_191 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_204 VDD gf180mcu_ocd_io__fill10x_204/one gf180mcu_ocd_io__fill10x_204/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_6 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_384 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_362 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_351 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_340 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_373 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__dvss_1 DVDD VSS VDD VSS gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_170 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_181 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_192 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_205 VDD gf180mcu_ocd_io__fill10x_205/one gf180mcu_ocd_io__fill10x_205/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_7 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_385 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_396 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_363 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_352 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_374 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_330 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__dvss_2 DVDD VSS VDD VSS gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_193 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_160 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_182 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_8 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_386 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_397 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_364 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_353 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_342 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_375 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_320 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_172 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_161 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_150 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_183 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_194 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__asig_5p0_0 DVDD VSS VDD analog_PAD[3] VSS gf180mcu_ocd_io__asig_5p0
Xgf180mcu_ocd_io__dvdd_1 VSS VDD VSS DVDD gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill5_9 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_398 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_387 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_365 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_354 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_343 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_376 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_332 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_321 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_162 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_173 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_140 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_151 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_184 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_195 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__asig_5p0_1 DVDD VSS VDD analog_PAD[2] VSS gf180mcu_ocd_io__asig_5p0
Xgf180mcu_ocd_io__in_s_0 DVDD gf180mcu_ocd_io__in_s_0/PD gf180mcu_ocd_io__in_s_0/PU
+ VDD gf180mcu_ocd_io__in_s_0/Y clk_PAD VSS VSS gf180mcu_ocd_io__in_s
Xgf180mcu_ocd_io__vss_0 DVDD VDD VSS VSS gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_388 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_399 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_366 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_344 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_377 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_322 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_333 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_311 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__dvss_5 DVDD VSS VDD VSS gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_130 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_174 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_141 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_152 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_185 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_196 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__asig_5p0_2 DVDD VSS VDD analog_PAD[0] VSS gf180mcu_ocd_io__asig_5p0
Xgf180mcu_ocd_io__cor_0 VDD DVDD VSS gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__dvdd_3 VSS VDD VSS DVDD gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_367 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_356 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_334 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_301 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_378 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_310x VDD gf180mcu_ocd_io__fill10_310x/one gf180mcu_ocd_io__fill10_310x/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_312 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_120 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_153 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_175 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_164 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_131 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_142 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_186 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__asig_5p0_3 DVDD VSS VDD analog_PAD[1] VSS gf180mcu_ocd_io__asig_5p0
Xgf180mcu_ocd_io__cor_1 VDD DVDD VSS gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__fill10x_190 VDD gf180mcu_ocd_io__fill10x_190/one gf180mcu_ocd_io__fill10x_190/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_368 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_346 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_357 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_335 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_302 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_379 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_324 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_313 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__dvss_7 DVDD VSS VDD VSS gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_110 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_165 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_132 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_143 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_198 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_176 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_187 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__vdd_0 DVDD VSS VDD VSS gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__cor_2 VDD DVDD VSS gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__dvdd_5 VSS VDD VSS DVDD gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10x_361 VDD gf180mcu_ocd_io__fill10x_361/one gf180mcu_ocd_io__fill10x_361/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_350 VDD gf180mcu_ocd_io__fill10x_350/one gf180mcu_ocd_io__fill10x_350/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__vss_3 DVDD VDD VSS VSS gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_369 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_358 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_347 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_303 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_325 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_314 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_199 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_111 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_133 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_166 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_155 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_122 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_144 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_188 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_100 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__cor_3 VDD DVDD VSS gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__dvdd_6 VSS VDD VSS DVDD gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10x_395 VDD gf180mcu_ocd_io__fill10x_395/one gf180mcu_ocd_io__fill10x_395/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__vss_4 DVDD VDD VSS VSS gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_359 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_348 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_337 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_304 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_326 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_315 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_101 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_112 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_167 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_156 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_178 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_123 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_134 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_145 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_189 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__vdd_2 DVDD VSS VDD VSS gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10x_341 VDD gf180mcu_ocd_io__fill10x_341/one gf180mcu_ocd_io__fill10x_341/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_171 VDD gf180mcu_ocd_io__fill10x_171/one gf180mcu_ocd_io__fill10x_171/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_349 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_338 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_305 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_327 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_316 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_168 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_157 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_135 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_124 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_146 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_179 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_331 VDD gf180mcu_ocd_io__fill10x_331/one gf180mcu_ocd_io__fill10x_331/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__vss_6 DVDD VDD VSS VSS gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_306 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_339 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_328 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_317 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_114 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_169 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_158 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_136 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_125 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_147 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__vdd_4 DVDD VSS VDD VSS gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10_90 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_329 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_104 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_115 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_159 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_137 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_148 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_355 VDD gf180mcu_ocd_io__fill10x_355/one gf180mcu_ocd_io__fill10x_355/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_300 VDD gf180mcu_ocd_io__fill10x_300/one gf180mcu_ocd_io__fill10x_300/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_91 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_80 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_163 VDD gf180mcu_ocd_io__fill10x_163/one gf180mcu_ocd_io__fill10x_163/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_319 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_308 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_116 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_105 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_127 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_149 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_345 VDD gf180mcu_ocd_io__fill10x_345/one gf180mcu_ocd_io__fill10x_345/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_323 VDD gf180mcu_ocd_io__fill10x_323/one gf180mcu_ocd_io__fill10x_323/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_92 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_70 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_81 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_389 VDD gf180mcu_ocd_io__fill10x_389/one gf180mcu_ocd_io__fill10x_389/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_197 VDD gf180mcu_ocd_io__fill10x_197/one gf180mcu_ocd_io__fill10x_197/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_309 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_117 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_139 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_128 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__vdd_7 DVDD VSS VDD VSS gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10_60 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_82 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_154 VDD gf180mcu_ocd_io__fill10x_154/one gf180mcu_ocd_io__fill10x_154/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_121 VDD gf180mcu_ocd_io__fill10x_121/one gf180mcu_ocd_io__fill10x_121/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_0 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_118 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_107 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_129 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_290 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_336 VDD gf180mcu_ocd_io__fill10x_336/one gf180mcu_ocd_io__fill10x_336/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_50 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_72 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_61 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_83 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_20 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10x_177 VDD gf180mcu_ocd_io__fill10x_177/one gf180mcu_ocd_io__fill10x_177/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_1 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_119 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_108 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_291 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_95 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_62 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_40 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_73 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_51 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_84 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_21 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill5_10 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_2 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_109 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_292 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_281 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_270 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_63 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_74 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_52 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_41 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_30 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_85 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_96 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_11 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10x_113 VDD gf180mcu_ocd_io__fill10x_113/one gf180mcu_ocd_io__fill10x_113/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_102 VDD gf180mcu_ocd_io__fill10x_102/one gf180mcu_ocd_io__fill10x_102/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_3 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_293 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_282 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_260 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_53 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_42 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_64 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_71 VDD gf180mcu_ocd_io__fill10x_71/one gf180mcu_ocd_io__fill10x_71/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_75 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_20 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_31 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_86 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_97 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_103 VDD gf180mcu_ocd_io__fill10x_103/one gf180mcu_ocd_io__fill10x_103/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_12 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_4 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_272 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_283 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_261 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_250 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_94 VDD gf180mcu_ocd_io__fill10x_94/one gf180mcu_ocd_io__fill10x_94/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_43 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_21 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_32 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_10 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_76 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_87 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_98 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_307 VDD gf180mcu_ocd_io__fill10x_307/one gf180mcu_ocd_io__fill10x_307/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_318 VDD gf180mcu_ocd_io__fill10x_318/one gf180mcu_ocd_io__fill10x_318/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_126 VDD gf180mcu_ocd_io__fill10x_126/one gf180mcu_ocd_io__fill10x_126/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_13 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_5 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_410 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_284 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_273 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_295 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_262 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_251 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_240 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_88 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_55 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_66 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_44 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_33 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_11 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_77 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_99 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_138 VDD gf180mcu_ocd_io__fill10x_138/one gf180mcu_ocd_io__fill10x_138/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill5_14 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_6 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_40 gf180mcu_ocd_io__bi_a_40/A gf180mcu_ocd_io__bi_a_40/ANA
+ gf180mcu_ocd_io__bi_a_40/CS DVDD gf180mcu_ocd_io__bi_a_40/IE gf180mcu_ocd_io__bi_a_40/OE
+ gf180mcu_ocd_io__bi_a_40/PD gf180mcu_ocd_io__bi_a_40/PDRV0 gf180mcu_ocd_io__bi_a_40/PDRV1
+ gf180mcu_ocd_io__bi_a_40/PU gf180mcu_ocd_io__bi_a_40/SL VDD gf180mcu_ocd_io__bi_a_40/Y
+ bidir_PAD[35] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_411 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_274 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_263 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_252 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_241 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_230 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_285 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_296 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_89 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_56 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_45 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_67 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_23 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_34 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_12 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_15 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10x_106 VDD gf180mcu_ocd_io__fill10x_106/one gf180mcu_ocd_io__fill10x_106/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_7 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_0 gf180mcu_ocd_io__bi_a_0/A gf180mcu_ocd_io__bi_a_0/ANA gf180mcu_ocd_io__bi_a_0/CS
+ DVDD gf180mcu_ocd_io__bi_a_0/IE gf180mcu_ocd_io__bi_a_0/OE gf180mcu_ocd_io__bi_a_0/PD
+ gf180mcu_ocd_io__bi_a_0/PDRV0 gf180mcu_ocd_io__bi_a_0/PDRV1 gf180mcu_ocd_io__bi_a_0/PU
+ gf180mcu_ocd_io__bi_a_0/SL VDD gf180mcu_ocd_io__bi_a_0/Y bidir_PAD[17] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_41 gf180mcu_ocd_io__bi_a_41/A gf180mcu_ocd_io__bi_a_41/ANA
+ gf180mcu_ocd_io__bi_a_41/CS DVDD gf180mcu_ocd_io__bi_a_41/IE gf180mcu_ocd_io__bi_a_41/OE
+ gf180mcu_ocd_io__bi_a_41/PD gf180mcu_ocd_io__bi_a_41/PDRV0 gf180mcu_ocd_io__bi_a_41/PDRV1
+ gf180mcu_ocd_io__bi_a_41/PU gf180mcu_ocd_io__bi_a_41/SL VDD gf180mcu_ocd_io__bi_a_41/Y
+ bidir_PAD[30] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_30 gf180mcu_ocd_io__bi_a_30/A gf180mcu_ocd_io__bi_a_30/ANA
+ gf180mcu_ocd_io__bi_a_30/CS DVDD gf180mcu_ocd_io__bi_a_30/IE gf180mcu_ocd_io__bi_a_30/OE
+ gf180mcu_ocd_io__bi_a_30/PD gf180mcu_ocd_io__bi_a_30/PDRV0 gf180mcu_ocd_io__bi_a_30/PDRV1
+ gf180mcu_ocd_io__bi_a_30/PU gf180mcu_ocd_io__bi_a_30/SL VDD gf180mcu_ocd_io__bi_a_30/Y
+ bidir_PAD[40] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_412 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_286 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_275 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_297 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_253 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_242 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_231 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_220 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_57 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_46 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_68 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_24 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_35 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_79 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_16 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_8 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_42 gf180mcu_ocd_io__bi_a_42/A gf180mcu_ocd_io__bi_a_42/ANA
+ gf180mcu_ocd_io__bi_a_42/CS DVDD gf180mcu_ocd_io__bi_a_42/IE gf180mcu_ocd_io__bi_a_42/OE
+ gf180mcu_ocd_io__bi_a_42/PD gf180mcu_ocd_io__bi_a_42/PDRV0 gf180mcu_ocd_io__bi_a_42/PDRV1
+ gf180mcu_ocd_io__bi_a_42/PU gf180mcu_ocd_io__bi_a_42/SL VDD gf180mcu_ocd_io__bi_a_42/Y
+ bidir_PAD[28] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_31 gf180mcu_ocd_io__bi_a_31/A gf180mcu_ocd_io__bi_a_31/ANA
+ gf180mcu_ocd_io__bi_a_31/CS DVDD gf180mcu_ocd_io__bi_a_31/IE gf180mcu_ocd_io__bi_a_31/OE
+ gf180mcu_ocd_io__bi_a_31/PD gf180mcu_ocd_io__bi_a_31/PDRV0 gf180mcu_ocd_io__bi_a_31/PDRV1
+ gf180mcu_ocd_io__bi_a_31/PU gf180mcu_ocd_io__bi_a_31/SL VDD gf180mcu_ocd_io__bi_a_31/Y
+ bidir_PAD[38] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_20 gf180mcu_ocd_io__bi_a_20/A gf180mcu_ocd_io__bi_a_20/ANA
+ gf180mcu_ocd_io__bi_a_20/CS DVDD gf180mcu_ocd_io__bi_a_20/IE gf180mcu_ocd_io__bi_a_20/OE
+ gf180mcu_ocd_io__bi_a_20/PD gf180mcu_ocd_io__bi_a_20/PDRV0 gf180mcu_ocd_io__bi_a_20/PDRV1
+ gf180mcu_ocd_io__bi_a_20/PU gf180mcu_ocd_io__bi_a_20/SL VDD gf180mcu_ocd_io__bi_a_20/Y
+ bidir_PAD[0] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_1 gf180mcu_ocd_io__bi_a_1/A gf180mcu_ocd_io__bi_a_1/ANA gf180mcu_ocd_io__bi_a_1/CS
+ DVDD gf180mcu_ocd_io__bi_a_1/IE gf180mcu_ocd_io__bi_a_1/OE gf180mcu_ocd_io__bi_a_1/PD
+ gf180mcu_ocd_io__bi_a_1/PDRV0 gf180mcu_ocd_io__bi_a_1/PDRV1 gf180mcu_ocd_io__bi_a_1/PU
+ gf180mcu_ocd_io__bi_a_1/SL VDD gf180mcu_ocd_io__bi_a_1/Y bidir_PAD[16] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_402 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_413 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_276 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_298 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_265 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_254 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_232 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_243 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_221 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_210 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_65 VDD gf180mcu_ocd_io__fill10x_65/one gf180mcu_ocd_io__fill10x_65/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_69 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_54 VDD gf180mcu_ocd_io__fill10x_54/one gf180mcu_ocd_io__fill10x_54/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_14 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_17 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_9 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_0 VDD gf180mcu_ocd_io__fill10x_0/one gf180mcu_ocd_io__fill10x_0/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__bi_a_43 gf180mcu_ocd_io__bi_a_43/A gf180mcu_ocd_io__bi_a_43/ANA
+ gf180mcu_ocd_io__bi_a_43/CS DVDD gf180mcu_ocd_io__bi_a_43/IE gf180mcu_ocd_io__bi_a_43/OE
+ gf180mcu_ocd_io__bi_a_43/PD gf180mcu_ocd_io__bi_a_43/PDRV0 gf180mcu_ocd_io__bi_a_43/PDRV1
+ gf180mcu_ocd_io__bi_a_43/PU gf180mcu_ocd_io__bi_a_43/SL VDD gf180mcu_ocd_io__bi_a_43/Y
+ bidir_PAD[27] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_32 gf180mcu_ocd_io__bi_a_32/A gf180mcu_ocd_io__bi_a_32/ANA
+ gf180mcu_ocd_io__bi_a_32/CS DVDD gf180mcu_ocd_io__bi_a_32/IE gf180mcu_ocd_io__bi_a_32/OE
+ gf180mcu_ocd_io__bi_a_32/PD gf180mcu_ocd_io__bi_a_32/PDRV0 gf180mcu_ocd_io__bi_a_32/PDRV1
+ gf180mcu_ocd_io__bi_a_32/PU gf180mcu_ocd_io__bi_a_32/SL VDD gf180mcu_ocd_io__bi_a_32/Y
+ bidir_PAD[23] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_21 gf180mcu_ocd_io__bi_a_21/A gf180mcu_ocd_io__bi_a_21/ANA
+ gf180mcu_ocd_io__bi_a_21/CS DVDD gf180mcu_ocd_io__bi_a_21/IE gf180mcu_ocd_io__bi_a_21/OE
+ gf180mcu_ocd_io__bi_a_21/PD gf180mcu_ocd_io__bi_a_21/PDRV0 gf180mcu_ocd_io__bi_a_21/PDRV1
+ gf180mcu_ocd_io__bi_a_21/PU gf180mcu_ocd_io__bi_a_21/SL VDD gf180mcu_ocd_io__bi_a_21/Y
+ bidir_PAD[1] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_2 gf180mcu_ocd_io__bi_a_2/A gf180mcu_ocd_io__bi_a_2/ANA gf180mcu_ocd_io__bi_a_2/CS
+ DVDD gf180mcu_ocd_io__bi_a_2/IE gf180mcu_ocd_io__bi_a_2/OE gf180mcu_ocd_io__bi_a_2/PD
+ gf180mcu_ocd_io__bi_a_2/PDRV0 gf180mcu_ocd_io__bi_a_2/PDRV1 gf180mcu_ocd_io__bi_a_2/PU
+ gf180mcu_ocd_io__bi_a_2/SL VDD gf180mcu_ocd_io__bi_a_2/Y bidir_PAD[15] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_10 gf180mcu_ocd_io__bi_a_10/A gf180mcu_ocd_io__bi_a_10/ANA
+ gf180mcu_ocd_io__bi_a_10/CS DVDD gf180mcu_ocd_io__bi_a_10/IE gf180mcu_ocd_io__bi_a_10/OE
+ gf180mcu_ocd_io__bi_a_10/PD gf180mcu_ocd_io__bi_a_10/PDRV0 gf180mcu_ocd_io__bi_a_10/PDRV1
+ gf180mcu_ocd_io__bi_a_10/PU gf180mcu_ocd_io__bi_a_10/SL VDD gf180mcu_ocd_io__bi_a_10/Y
+ bidir_PAD[19] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_280 VDD gf180mcu_ocd_io__fill10x_280/one gf180mcu_ocd_io__fill10x_280/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_403 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_288 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_277 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_299 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_255 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_244 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_233 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_222 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_211 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_200 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_48 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_26 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_22 VDD gf180mcu_ocd_io__fill10x_22/one gf180mcu_ocd_io__fill10x_22/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_15 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_37 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_18 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__bi_a_44 gf180mcu_ocd_io__bi_a_44/A gf180mcu_ocd_io__bi_a_44/ANA
+ gf180mcu_ocd_io__bi_a_44/CS DVDD gf180mcu_ocd_io__bi_a_44/IE gf180mcu_ocd_io__bi_a_44/OE
+ gf180mcu_ocd_io__bi_a_44/PD gf180mcu_ocd_io__bi_a_44/PDRV0 gf180mcu_ocd_io__bi_a_44/PDRV1
+ gf180mcu_ocd_io__bi_a_44/PU gf180mcu_ocd_io__bi_a_44/SL VDD gf180mcu_ocd_io__bi_a_44/Y
+ bidir_PAD[26] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_22 gf180mcu_ocd_io__bi_a_22/A gf180mcu_ocd_io__bi_a_22/ANA
+ gf180mcu_ocd_io__bi_a_22/CS DVDD gf180mcu_ocd_io__bi_a_22/IE gf180mcu_ocd_io__bi_a_22/OE
+ gf180mcu_ocd_io__bi_a_22/PD gf180mcu_ocd_io__bi_a_22/PDRV0 gf180mcu_ocd_io__bi_a_22/PDRV1
+ gf180mcu_ocd_io__bi_a_22/PU gf180mcu_ocd_io__bi_a_22/SL VDD gf180mcu_ocd_io__bi_a_22/Y
+ bidir_PAD[45] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_33 gf180mcu_ocd_io__bi_a_33/A gf180mcu_ocd_io__bi_a_33/ANA
+ gf180mcu_ocd_io__bi_a_33/CS DVDD gf180mcu_ocd_io__bi_a_33/IE gf180mcu_ocd_io__bi_a_33/OE
+ gf180mcu_ocd_io__bi_a_33/PD gf180mcu_ocd_io__bi_a_33/PDRV0 gf180mcu_ocd_io__bi_a_33/PDRV1
+ gf180mcu_ocd_io__bi_a_33/PU gf180mcu_ocd_io__bi_a_33/SL VDD gf180mcu_ocd_io__bi_a_33/Y
+ bidir_PAD[22] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_3 gf180mcu_ocd_io__bi_a_3/A gf180mcu_ocd_io__bi_a_3/ANA gf180mcu_ocd_io__bi_a_3/CS
+ DVDD gf180mcu_ocd_io__bi_a_3/IE gf180mcu_ocd_io__bi_a_3/OE gf180mcu_ocd_io__bi_a_3/PD
+ gf180mcu_ocd_io__bi_a_3/PDRV0 gf180mcu_ocd_io__bi_a_3/PDRV1 gf180mcu_ocd_io__bi_a_3/PU
+ gf180mcu_ocd_io__bi_a_3/SL VDD gf180mcu_ocd_io__bi_a_3/Y bidir_PAD[14] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_11 gf180mcu_ocd_io__bi_a_11/A gf180mcu_ocd_io__bi_a_11/ANA
+ gf180mcu_ocd_io__bi_a_11/CS DVDD gf180mcu_ocd_io__bi_a_11/IE gf180mcu_ocd_io__bi_a_11/OE
+ gf180mcu_ocd_io__bi_a_11/PD gf180mcu_ocd_io__bi_a_11/PDRV0 gf180mcu_ocd_io__bi_a_11/PDRV1
+ gf180mcu_ocd_io__bi_a_11/PU gf180mcu_ocd_io__bi_a_11/SL VDD gf180mcu_ocd_io__bi_a_11/Y
+ bidir_PAD[18] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_404 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_289 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_278 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_256 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_245 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_267 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_234 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_223 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_212 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_201 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_78 VDD gf180mcu_ocd_io__fill10x_78/one gf180mcu_ocd_io__fill10x_78/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_49 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_27 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_16 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_38 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_19 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__bi_a_45 gf180mcu_ocd_io__bi_a_45/A gf180mcu_ocd_io__bi_a_45/ANA
+ gf180mcu_ocd_io__bi_a_45/CS DVDD gf180mcu_ocd_io__bi_a_45/IE gf180mcu_ocd_io__bi_a_45/OE
+ gf180mcu_ocd_io__bi_a_45/PD gf180mcu_ocd_io__bi_a_45/PDRV0 gf180mcu_ocd_io__bi_a_45/PDRV1
+ gf180mcu_ocd_io__bi_a_45/PU gf180mcu_ocd_io__bi_a_45/SL VDD gf180mcu_ocd_io__bi_a_45/Y
+ bidir_PAD[29] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_23 gf180mcu_ocd_io__bi_a_23/A gf180mcu_ocd_io__bi_a_23/ANA
+ gf180mcu_ocd_io__bi_a_23/CS DVDD gf180mcu_ocd_io__bi_a_23/IE gf180mcu_ocd_io__bi_a_23/OE
+ gf180mcu_ocd_io__bi_a_23/PD gf180mcu_ocd_io__bi_a_23/PDRV0 gf180mcu_ocd_io__bi_a_23/PDRV1
+ gf180mcu_ocd_io__bi_a_23/PU gf180mcu_ocd_io__bi_a_23/SL VDD gf180mcu_ocd_io__bi_a_23/Y
+ bidir_PAD[43] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_34 gf180mcu_ocd_io__bi_a_34/A gf180mcu_ocd_io__bi_a_34/ANA
+ gf180mcu_ocd_io__bi_a_34/CS DVDD gf180mcu_ocd_io__bi_a_34/IE gf180mcu_ocd_io__bi_a_34/OE
+ gf180mcu_ocd_io__bi_a_34/PD gf180mcu_ocd_io__bi_a_34/PDRV0 gf180mcu_ocd_io__bi_a_34/PDRV1
+ gf180mcu_ocd_io__bi_a_34/PU gf180mcu_ocd_io__bi_a_34/SL VDD gf180mcu_ocd_io__bi_a_34/Y
+ bidir_PAD[24] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_12 gf180mcu_ocd_io__bi_a_12/A gf180mcu_ocd_io__bi_a_12/ANA
+ gf180mcu_ocd_io__bi_a_12/CS DVDD gf180mcu_ocd_io__bi_a_12/IE gf180mcu_ocd_io__bi_a_12/OE
+ gf180mcu_ocd_io__bi_a_12/PD gf180mcu_ocd_io__bi_a_12/PDRV0 gf180mcu_ocd_io__bi_a_12/PDRV1
+ gf180mcu_ocd_io__bi_a_12/PU gf180mcu_ocd_io__bi_a_12/SL VDD gf180mcu_ocd_io__bi_a_12/Y
+ bidir_PAD[20] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_4 gf180mcu_ocd_io__bi_a_4/A gf180mcu_ocd_io__bi_a_4/ANA gf180mcu_ocd_io__bi_a_4/CS
+ DVDD gf180mcu_ocd_io__bi_a_4/IE gf180mcu_ocd_io__bi_a_4/OE gf180mcu_ocd_io__bi_a_4/PD
+ gf180mcu_ocd_io__bi_a_4/PDRV0 gf180mcu_ocd_io__bi_a_4/PDRV1 gf180mcu_ocd_io__bi_a_4/PU
+ gf180mcu_ocd_io__bi_a_4/SL VDD gf180mcu_ocd_io__bi_a_4/Y bidir_PAD[10] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_271 VDD gf180mcu_ocd_io__fill10x_271/one gf180mcu_ocd_io__fill10x_271/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_405 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_279 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_257 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_246 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_268 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_235 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_224 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_213 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_202 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_13 VDD gf180mcu_ocd_io__fill10x_13/one gf180mcu_ocd_io__fill10x_13/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_39 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_28 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_17 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_24 gf180mcu_ocd_io__bi_a_24/A gf180mcu_ocd_io__bi_a_24/ANA
+ gf180mcu_ocd_io__bi_a_24/CS DVDD gf180mcu_ocd_io__bi_a_24/IE gf180mcu_ocd_io__bi_a_24/OE
+ gf180mcu_ocd_io__bi_a_24/PD gf180mcu_ocd_io__bi_a_24/PDRV0 gf180mcu_ocd_io__bi_a_24/PDRV1
+ gf180mcu_ocd_io__bi_a_24/PU gf180mcu_ocd_io__bi_a_24/SL VDD gf180mcu_ocd_io__bi_a_24/Y
+ bidir_PAD[42] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_35 gf180mcu_ocd_io__bi_a_35/A gf180mcu_ocd_io__bi_a_35/ANA
+ gf180mcu_ocd_io__bi_a_35/CS DVDD gf180mcu_ocd_io__bi_a_35/IE gf180mcu_ocd_io__bi_a_35/OE
+ gf180mcu_ocd_io__bi_a_35/PD gf180mcu_ocd_io__bi_a_35/PDRV0 gf180mcu_ocd_io__bi_a_35/PDRV1
+ gf180mcu_ocd_io__bi_a_35/PU gf180mcu_ocd_io__bi_a_35/SL VDD gf180mcu_ocd_io__bi_a_35/Y
+ bidir_PAD[25] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_13 gf180mcu_ocd_io__bi_a_13/A gf180mcu_ocd_io__bi_a_13/ANA
+ gf180mcu_ocd_io__bi_a_13/CS DVDD gf180mcu_ocd_io__bi_a_13/IE gf180mcu_ocd_io__bi_a_13/OE
+ gf180mcu_ocd_io__bi_a_13/PD gf180mcu_ocd_io__bi_a_13/PDRV0 gf180mcu_ocd_io__bi_a_13/PDRV1
+ gf180mcu_ocd_io__bi_a_13/PU gf180mcu_ocd_io__bi_a_13/SL VDD gf180mcu_ocd_io__bi_a_13/Y
+ bidir_PAD[21] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_5 gf180mcu_ocd_io__bi_a_5/A gf180mcu_ocd_io__bi_a_5/ANA gf180mcu_ocd_io__bi_a_5/CS
+ DVDD gf180mcu_ocd_io__bi_a_5/IE gf180mcu_ocd_io__bi_a_5/OE gf180mcu_ocd_io__bi_a_5/PD
+ gf180mcu_ocd_io__bi_a_5/PDRV0 gf180mcu_ocd_io__bi_a_5/PDRV1 gf180mcu_ocd_io__bi_a_5/PU
+ gf180mcu_ocd_io__bi_a_5/SL VDD gf180mcu_ocd_io__bi_a_5/Y bidir_PAD[8] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_294 VDD gf180mcu_ocd_io__fill10x_294/one gf180mcu_ocd_io__fill10x_294/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_406 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_25 VDD gf180mcu_ocd_io__fill10x_25/one gf180mcu_ocd_io__fill10x_25/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_36 VDD gf180mcu_ocd_io__fill10x_36/one gf180mcu_ocd_io__fill10x_36/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_269 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_236 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_225 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_214 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_203 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_58 VDD gf180mcu_ocd_io__fill10x_58/one gf180mcu_ocd_io__fill10x_58/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_47 VDD gf180mcu_ocd_io__fill10x_47/one gf180mcu_ocd_io__fill10x_47/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_18 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_29 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_6 gf180mcu_ocd_io__bi_a_6/A gf180mcu_ocd_io__bi_a_6/ANA gf180mcu_ocd_io__bi_a_6/CS
+ DVDD gf180mcu_ocd_io__bi_a_6/IE gf180mcu_ocd_io__bi_a_6/OE gf180mcu_ocd_io__bi_a_6/PD
+ gf180mcu_ocd_io__bi_a_6/PDRV0 gf180mcu_ocd_io__bi_a_6/PDRV1 gf180mcu_ocd_io__bi_a_6/PU
+ gf180mcu_ocd_io__bi_a_6/SL VDD gf180mcu_ocd_io__bi_a_6/Y bidir_PAD[11] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_36 gf180mcu_ocd_io__bi_a_36/A gf180mcu_ocd_io__bi_a_36/ANA
+ gf180mcu_ocd_io__bi_a_36/CS DVDD gf180mcu_ocd_io__bi_a_36/IE gf180mcu_ocd_io__bi_a_36/OE
+ gf180mcu_ocd_io__bi_a_36/PD gf180mcu_ocd_io__bi_a_36/PDRV0 gf180mcu_ocd_io__bi_a_36/PDRV1
+ gf180mcu_ocd_io__bi_a_36/PU gf180mcu_ocd_io__bi_a_36/SL VDD gf180mcu_ocd_io__bi_a_36/Y
+ bidir_PAD[31] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_25 gf180mcu_ocd_io__bi_a_25/A gf180mcu_ocd_io__bi_a_25/ANA
+ gf180mcu_ocd_io__bi_a_25/CS DVDD gf180mcu_ocd_io__bi_a_25/IE gf180mcu_ocd_io__bi_a_25/OE
+ gf180mcu_ocd_io__bi_a_25/PD gf180mcu_ocd_io__bi_a_25/PDRV0 gf180mcu_ocd_io__bi_a_25/PDRV1
+ gf180mcu_ocd_io__bi_a_25/PU gf180mcu_ocd_io__bi_a_25/SL VDD gf180mcu_ocd_io__bi_a_25/Y
+ bidir_PAD[44] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_14 gf180mcu_ocd_io__bi_a_14/A gf180mcu_ocd_io__bi_a_14/ANA
+ gf180mcu_ocd_io__bi_a_14/CS DVDD gf180mcu_ocd_io__bi_a_14/IE gf180mcu_ocd_io__bi_a_14/OE
+ gf180mcu_ocd_io__bi_a_14/PD gf180mcu_ocd_io__bi_a_14/PDRV0 gf180mcu_ocd_io__bi_a_14/PDRV1
+ gf180mcu_ocd_io__bi_a_14/PU gf180mcu_ocd_io__bi_a_14/SL VDD gf180mcu_ocd_io__bi_a_14/Y
+ bidir_PAD[3] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_407 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_259 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_248 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_237 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_226 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_215 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_59 VDD gf180mcu_ocd_io__fill10x_59/one gf180mcu_ocd_io__fill10x_59/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_19 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_400 VDD gf180mcu_ocd_io__fill10x_400/one gf180mcu_ocd_io__fill10x_400/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__bi_a_37 gf180mcu_ocd_io__bi_a_37/A gf180mcu_ocd_io__bi_a_37/ANA
+ gf180mcu_ocd_io__bi_a_37/CS DVDD gf180mcu_ocd_io__bi_a_37/IE gf180mcu_ocd_io__bi_a_37/OE
+ gf180mcu_ocd_io__bi_a_37/PD gf180mcu_ocd_io__bi_a_37/PDRV0 gf180mcu_ocd_io__bi_a_37/PDRV1
+ gf180mcu_ocd_io__bi_a_37/PU gf180mcu_ocd_io__bi_a_37/SL VDD gf180mcu_ocd_io__bi_a_37/Y
+ bidir_PAD[32] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_26 gf180mcu_ocd_io__bi_a_26/A gf180mcu_ocd_io__bi_a_26/ANA
+ gf180mcu_ocd_io__bi_a_26/CS DVDD gf180mcu_ocd_io__bi_a_26/IE gf180mcu_ocd_io__bi_a_26/OE
+ gf180mcu_ocd_io__bi_a_26/PD gf180mcu_ocd_io__bi_a_26/PDRV0 gf180mcu_ocd_io__bi_a_26/PDRV1
+ gf180mcu_ocd_io__bi_a_26/PU gf180mcu_ocd_io__bi_a_26/SL VDD gf180mcu_ocd_io__bi_a_26/Y
+ bidir_PAD[36] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_15 gf180mcu_ocd_io__bi_a_15/A gf180mcu_ocd_io__bi_a_15/ANA
+ gf180mcu_ocd_io__bi_a_15/CS DVDD gf180mcu_ocd_io__bi_a_15/IE gf180mcu_ocd_io__bi_a_15/OE
+ gf180mcu_ocd_io__bi_a_15/PD gf180mcu_ocd_io__bi_a_15/PDRV0 gf180mcu_ocd_io__bi_a_15/PDRV1
+ gf180mcu_ocd_io__bi_a_15/PU gf180mcu_ocd_io__bi_a_15/SL VDD gf180mcu_ocd_io__bi_a_15/Y
+ bidir_PAD[6] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_7 gf180mcu_ocd_io__bi_a_7/A gf180mcu_ocd_io__bi_a_7/ANA gf180mcu_ocd_io__bi_a_7/CS
+ DVDD gf180mcu_ocd_io__bi_a_7/IE gf180mcu_ocd_io__bi_a_7/OE gf180mcu_ocd_io__bi_a_7/PD
+ gf180mcu_ocd_io__bi_a_7/PDRV0 gf180mcu_ocd_io__bi_a_7/PDRV1 gf180mcu_ocd_io__bi_a_7/PU
+ gf180mcu_ocd_io__bi_a_7/SL VDD gf180mcu_ocd_io__bi_a_7/Y bidir_PAD[13] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_408 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_249 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_238 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_227 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_216 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__in_c_0 DVDD gf180mcu_ocd_io__in_c_0/PD gf180mcu_ocd_io__in_c_0/PU
+ VDD gf180mcu_ocd_io__in_c_0/Y rst_n_PAD VSS VSS gf180mcu_ocd_io__in_c
Xgf180mcu_ocd_io__fill10x_401 VDD gf180mcu_ocd_io__fill10x_401/one gf180mcu_ocd_io__fill10x_401/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__bi_a_38 gf180mcu_ocd_io__bi_a_38/A gf180mcu_ocd_io__bi_a_38/ANA
+ gf180mcu_ocd_io__bi_a_38/CS DVDD gf180mcu_ocd_io__bi_a_38/IE gf180mcu_ocd_io__bi_a_38/OE
+ gf180mcu_ocd_io__bi_a_38/PD gf180mcu_ocd_io__bi_a_38/PDRV0 gf180mcu_ocd_io__bi_a_38/PDRV1
+ gf180mcu_ocd_io__bi_a_38/PU gf180mcu_ocd_io__bi_a_38/SL VDD gf180mcu_ocd_io__bi_a_38/Y
+ bidir_PAD[34] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_27 gf180mcu_ocd_io__bi_a_27/A gf180mcu_ocd_io__bi_a_27/ANA
+ gf180mcu_ocd_io__bi_a_27/CS DVDD gf180mcu_ocd_io__bi_a_27/IE gf180mcu_ocd_io__bi_a_27/OE
+ gf180mcu_ocd_io__bi_a_27/PD gf180mcu_ocd_io__bi_a_27/PDRV0 gf180mcu_ocd_io__bi_a_27/PDRV1
+ gf180mcu_ocd_io__bi_a_27/PU gf180mcu_ocd_io__bi_a_27/SL VDD gf180mcu_ocd_io__bi_a_27/Y
+ bidir_PAD[39] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_16 gf180mcu_ocd_io__bi_a_16/A gf180mcu_ocd_io__bi_a_16/ANA
+ gf180mcu_ocd_io__bi_a_16/CS DVDD gf180mcu_ocd_io__bi_a_16/IE gf180mcu_ocd_io__bi_a_16/OE
+ gf180mcu_ocd_io__bi_a_16/PD gf180mcu_ocd_io__bi_a_16/PDRV0 gf180mcu_ocd_io__bi_a_16/PDRV1
+ gf180mcu_ocd_io__bi_a_16/PU gf180mcu_ocd_io__bi_a_16/SL VDD gf180mcu_ocd_io__bi_a_16/Y
+ bidir_PAD[7] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_8 gf180mcu_ocd_io__bi_a_8/A gf180mcu_ocd_io__bi_a_8/ANA gf180mcu_ocd_io__bi_a_8/CS
+ DVDD gf180mcu_ocd_io__bi_a_8/IE gf180mcu_ocd_io__bi_a_8/OE gf180mcu_ocd_io__bi_a_8/PD
+ gf180mcu_ocd_io__bi_a_8/PDRV0 gf180mcu_ocd_io__bi_a_8/PDRV1 gf180mcu_ocd_io__bi_a_8/PU
+ gf180mcu_ocd_io__bi_a_8/SL VDD gf180mcu_ocd_io__bi_a_8/Y bidir_PAD[12] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_264 VDD gf180mcu_ocd_io__fill10x_264/one gf180mcu_ocd_io__fill10x_264/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_409 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_239 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_228 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_217 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_206 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_0 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__in_c_1 DVDD gf180mcu_ocd_io__in_c_1/PD gf180mcu_ocd_io__in_c_1/PU
+ VDD gf180mcu_ocd_io__in_c_1/Y input_PAD[3] VSS VSS gf180mcu_ocd_io__in_c
Xgf180mcu_ocd_io__bi_a_39 gf180mcu_ocd_io__bi_a_39/A gf180mcu_ocd_io__bi_a_39/ANA
+ gf180mcu_ocd_io__bi_a_39/CS DVDD gf180mcu_ocd_io__bi_a_39/IE gf180mcu_ocd_io__bi_a_39/OE
+ gf180mcu_ocd_io__bi_a_39/PD gf180mcu_ocd_io__bi_a_39/PDRV0 gf180mcu_ocd_io__bi_a_39/PDRV1
+ gf180mcu_ocd_io__bi_a_39/PU gf180mcu_ocd_io__bi_a_39/SL VDD gf180mcu_ocd_io__bi_a_39/Y
+ bidir_PAD[33] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_28 gf180mcu_ocd_io__bi_a_28/A gf180mcu_ocd_io__bi_a_28/ANA
+ gf180mcu_ocd_io__bi_a_28/CS DVDD gf180mcu_ocd_io__bi_a_28/IE gf180mcu_ocd_io__bi_a_28/OE
+ gf180mcu_ocd_io__bi_a_28/PD gf180mcu_ocd_io__bi_a_28/PDRV0 gf180mcu_ocd_io__bi_a_28/PDRV1
+ gf180mcu_ocd_io__bi_a_28/PU gf180mcu_ocd_io__bi_a_28/SL VDD gf180mcu_ocd_io__bi_a_28/Y
+ bidir_PAD[37] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_17 gf180mcu_ocd_io__bi_a_17/A gf180mcu_ocd_io__bi_a_17/ANA
+ gf180mcu_ocd_io__bi_a_17/CS DVDD gf180mcu_ocd_io__bi_a_17/IE gf180mcu_ocd_io__bi_a_17/OE
+ gf180mcu_ocd_io__bi_a_17/PD gf180mcu_ocd_io__bi_a_17/PDRV0 gf180mcu_ocd_io__bi_a_17/PDRV1
+ gf180mcu_ocd_io__bi_a_17/PU gf180mcu_ocd_io__bi_a_17/SL VDD gf180mcu_ocd_io__bi_a_17/Y
+ bidir_PAD[4] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_9 gf180mcu_ocd_io__bi_a_9/A gf180mcu_ocd_io__bi_a_9/ANA gf180mcu_ocd_io__bi_a_9/CS
+ DVDD gf180mcu_ocd_io__bi_a_9/IE gf180mcu_ocd_io__bi_a_9/OE gf180mcu_ocd_io__bi_a_9/PD
+ gf180mcu_ocd_io__bi_a_9/PDRV0 gf180mcu_ocd_io__bi_a_9/PDRV1 gf180mcu_ocd_io__bi_a_9/PU
+ gf180mcu_ocd_io__bi_a_9/SL VDD gf180mcu_ocd_io__bi_a_9/Y bidir_PAD[9] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_287 VDD gf180mcu_ocd_io__fill10x_287/one gf180mcu_ocd_io__fill10x_287/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_229 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_218 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_207 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_1 VDD VSS DVDD VSS gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__in_c_2 DVDD gf180mcu_ocd_io__in_c_2/PD gf180mcu_ocd_io__in_c_2/PU
+ VDD gf180mcu_ocd_io__in_c_2/Y input_PAD[2] VSS VSS gf180mcu_ocd_io__in_c
Xgf180mcu_ocd_io__fill10_390 VDD VSS DVDD VSS gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_29 gf180mcu_ocd_io__bi_a_29/A gf180mcu_ocd_io__bi_a_29/ANA
+ gf180mcu_ocd_io__bi_a_29/CS DVDD gf180mcu_ocd_io__bi_a_29/IE gf180mcu_ocd_io__bi_a_29/OE
+ gf180mcu_ocd_io__bi_a_29/PD gf180mcu_ocd_io__bi_a_29/PDRV0 gf180mcu_ocd_io__bi_a_29/PDRV1
+ gf180mcu_ocd_io__bi_a_29/PU gf180mcu_ocd_io__bi_a_29/SL VDD gf180mcu_ocd_io__bi_a_29/Y
+ bidir_PAD[41] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__bi_a_18 gf180mcu_ocd_io__bi_a_18/A gf180mcu_ocd_io__bi_a_18/ANA
+ gf180mcu_ocd_io__bi_a_18/CS DVDD gf180mcu_ocd_io__bi_a_18/IE gf180mcu_ocd_io__bi_a_18/OE
+ gf180mcu_ocd_io__bi_a_18/PD gf180mcu_ocd_io__bi_a_18/PDRV0 gf180mcu_ocd_io__bi_a_18/PDRV1
+ gf180mcu_ocd_io__bi_a_18/PU gf180mcu_ocd_io__bi_a_18/SL VDD gf180mcu_ocd_io__bi_a_18/Y
+ bidir_PAD[5] VSS VSS gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_266 VDD gf180mcu_ocd_io__fill10x_266/one gf180mcu_ocd_io__fill10x_266/zero
+ DVDD VSS VSS gf180mcu_ocd_io__fill10x
.ends

.subckt gf180mcu_ocd_sram_test
Xgf180mcu_ocd_ip_sram__sram512x8m8wm1_0 GWEN Q7_512_2 Q6_512_2 Q5_512_2 Q4_512_2 Q3_512_2
+ Q2_512_2 Q1_512_2 D6 WEN7 WEN6 WEN5 WEN4 WEN3 A0 D1 A1 A2 D3 A3 A4 D5 A5 A6 D7 A7
+ A8 ENA_512_2 VSS WEN0 CLK WEN1 WEN2 Q0_512_2 gf180mcu_ocd_ip_sram__sram512x8m8wm1
Xgf180mcu_ocd_ip_sram__sram512x8m8wm1_1 GWEN Q7_512_1 Q6_512_1 Q5_512_1 Q4_512_1 Q3_512_1
+ Q2_512_1 Q1_512_1 D6 WEN7 WEN6 WEN5 WEN4 WEN3 A0 D1 A1 A2 D3 A3 A4 D5 A5 A6 D7 A7
+ A8 ENA_512_1 VSS WEN0 CLK WEN1 WEN2 Q0_512_1 gf180mcu_ocd_ip_sram__sram512x8m8wm1
Xlvlshift_down_0 D6 simple_por_0/VDD simple_por_0/por VSS lvlshift_down_0/YL lvlshift_down
Xsimple_por_0 simple_por_0/VDD simple_por_0/porb simple_por_0/por VSS simple_por
Xgf180mcu_ocd_ip_sram__sram256x8m8wm1_0 A7 A6 A5 A4 A3 A2 A1 A0 ENA_256_1 CLK D7 D5
+ D3 D1 GWEN Q7_256_1 Q6_256_1 Q5_256_1 Q4_256_1 Q3_256_1 Q2_256_1 Q1_256_1 Q0_256_1
+ D6 WEN7 WEN6 WEN5 WEN4 WEN3 WEN2 WEN1 WEN0 VSS gf180mcu_ocd_ip_sram__sram256x8m8wm1
Xgf180mcu_ocd_ip_sram__sram256x8m8wm1_1 A7 A6 A5 A4 A3 A2 A1 A0 ENA_256_2 CLK D7 D5
+ D3 D1 GWEN Q7_256_2 Q6_256_2 Q5_256_2 Q4_256_2 Q3_256_2 Q2_256_2 Q1_256_2 Q0_256_2
+ D6 WEN7 WEN6 WEN5 WEN4 WEN3 WEN2 WEN1 WEN0 VSS gf180mcu_ocd_ip_sram__sram256x8m8wm1
Xocd_mux_array_0 select_256 Q0_256_1 Q1_256_1 Q2_256_1 Q3_256_1 Q4_256_1 Q5_256_1
+ Q6_256_1 Q7_256_1 Q0_256_2 Q1_256_2 Q2_256_2 Q3_256_2 Q4_256_2 Q5_256_2 Q6_256_2
+ Q7_256_2 ocd_mux_array_0/Y[7] ocd_mux_array_0/Y[3] ocd_mux_array_0/Y[5] ocd_mux_array_0/Y[1]
+ ocd_mux_array_0/Y[6] D6 ocd_mux_array_0/Y[4] ocd_mux_array_0/Y[0] VSS ocd_mux_array_0/Y[2]
+ ocd_mux_array
Xocd_mux_array_1 select_512 Q0_512_1 Q1_512_1 Q2_512_1 Q3_512_1 Q4_512_1 Q5_512_1
+ Q6_512_1 Q7_512_1 Q0_512_2 Q1_512_2 Q2_512_2 Q3_512_2 Q4_512_2 Q5_512_2 Q6_512_2
+ Q7_512_2 ocd_mux_array_1/Y[7] ocd_mux_array_1/Y[3] ocd_mux_array_1/Y[5] ocd_mux_array_1/Y[1]
+ ocd_mux_array_1/Y[6] D6 ocd_mux_array_1/Y[4] ocd_mux_array_1/Y[0] VSS ocd_mux_array_1/Y[2]
+ ocd_mux_array
Xchip_half_frame_0 simple_por_0/VDD chip_half_frame_0/analog_PAD[0] chip_half_frame_0/analog_PAD[1]
+ chip_half_frame_0/analog_PAD[2] chip_half_frame_0/analog_PAD[3] chip_half_frame_0/input_PAD[0]
+ chip_half_frame_0/input_PAD[1] chip_half_frame_0/input_PAD[2] chip_half_frame_0/input_PAD[3]
+ chip_half_frame_0/clk_PAD chip_half_frame_0/rst_n_PAD chip_half_frame_0/bidir_PAD[0]
+ chip_half_frame_0/bidir_PAD[1] chip_half_frame_0/bidir_PAD[2] chip_half_frame_0/bidir_PAD[3]
+ chip_half_frame_0/bidir_PAD[4] chip_half_frame_0/bidir_PAD[5] chip_half_frame_0/bidir_PAD[6]
+ chip_half_frame_0/bidir_PAD[7] chip_half_frame_0/bidir_PAD[8] chip_half_frame_0/bidir_PAD[9]
+ chip_half_frame_0/bidir_PAD[10] chip_half_frame_0/bidir_PAD[11] chip_half_frame_0/bidir_PAD[12]
+ chip_half_frame_0/bidir_PAD[13] chip_half_frame_0/bidir_PAD[14] chip_half_frame_0/bidir_PAD[15]
+ chip_half_frame_0/bidir_PAD[16] chip_half_frame_0/bidir_PAD[17] chip_half_frame_0/bidir_PAD[18]
+ chip_half_frame_0/bidir_PAD[19] chip_half_frame_0/bidir_PAD[20] chip_half_frame_0/bidir_PAD[21]
+ chip_half_frame_0/bidir_PAD[22] chip_half_frame_0/bidir_PAD[23] chip_half_frame_0/bidir_PAD[24]
+ chip_half_frame_0/bidir_PAD[25] chip_half_frame_0/bidir_PAD[26] chip_half_frame_0/bidir_PAD[27]
+ chip_half_frame_0/bidir_PAD[28] chip_half_frame_0/bidir_PAD[29] chip_half_frame_0/bidir_PAD[30]
+ chip_half_frame_0/bidir_PAD[31] chip_half_frame_0/bidir_PAD[32] chip_half_frame_0/bidir_PAD[33]
+ chip_half_frame_0/bidir_PAD[34] chip_half_frame_0/bidir_PAD[35] chip_half_frame_0/bidir_PAD[36]
+ chip_half_frame_0/bidir_PAD[37] chip_half_frame_0/bidir_PAD[38] chip_half_frame_0/bidir_PAD[39]
+ chip_half_frame_0/bidir_PAD[40] chip_half_frame_0/bidir_PAD[41] chip_half_frame_0/bidir_PAD[42]
+ chip_half_frame_0/bidir_PAD[43] chip_half_frame_0/bidir_PAD[44] chip_half_frame_0/bidir_PAD[45]
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/IE
+ ENA_512_1 D1 chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/OE
+ WEN6 A5 chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A
+ select_256 chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_1/PD chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A ENA_256_2 chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/OE
+ WEN5 chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL ocd_mux_array_0/Y[1] chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A D6 CLK A2 chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/OE
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_0/PU select_512 chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL
+ ocd_mux_array_0/Y[4] chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL chip_half_frame_0/gf180mcu_ocd_io__in_c_3/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A chip_half_frame_0/gf180mcu_ocd_io__in_c_0/Y
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A
+ D3 chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A
+ ocd_mux_array_1/Y[0] chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/IE
+ A7 chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A
+ ocd_mux_array_0/Y[7] chip_half_frame_0/gf180mcu_ocd_io__in_c_3/PU chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL
+ D6 chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/IE chip_half_frame_0/gf180mcu_ocd_io__in_c_2/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/IE WEN0 chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A
+ ocd_mux_array_1/Y[5] chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A
+ WEN7 A4 chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL A8 chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL chip_half_frame_0/gf180mcu_ocd_io__in_c_1/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A
+ ocd_mux_array_1/Y[2] chip_half_frame_0/gf180mcu_ocd_io__in_c_0/PU chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/IE
+ ENA_512_2 chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/IE chip_half_frame_0/gf180mcu_ocd_io__in_s_0/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL ocd_mux_array_0/Y[2] chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A WEN3 chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/OE
+ ocd_mux_array_1/Y[6] chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/IE D5 chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/OE A1 chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_1/PD chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL ENA_256_1 chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/OE
+ GWEN chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/IE
+ chip_half_frame_0/gf180mcu_ocd_io__in_s_0/PU chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ ocd_mux_array_0/Y[5] chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_0/PD chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_1/PU chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A D6 chip_half_frame_0/gf180mcu_ocd_io__in_s_0/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/OE
+ ocd_mux_array_1/Y[1] chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__in_c_2/PU
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/OE ocd_mux_array_1/Y[3] chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ A6 chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_2/PU WEN4 chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ ocd_mux_array_0/Y[0] chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_15/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_6/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL chip_half_frame_0/gf180mcu_ocd_io__in_c_0/PD
+ D7 chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A
+ A3 chip_half_frame_0/gf180mcu_ocd_io__bi_a_5/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_8/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_45/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_7/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_37/SL
+ ocd_mux_array_0/Y[3] chip_half_frame_0/gf180mcu_ocd_io__bi_a_42/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/OE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_9/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_39/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/SL
+ WEN1 chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_34/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_2/A
+ chip_half_frame_0/gf180mcu_ocd_io__in_c_3/PU chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A
+ ocd_mux_array_1/Y[7] chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_18/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL D6 chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_26/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_36/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_20/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_31/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_29/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ D6 chip_half_frame_0/gf180mcu_ocd_io__bi_a_28/SL lvlshift_down_0/YL chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_23/SL A0 chip_half_frame_0/gf180mcu_ocd_io__bi_a_33/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_21/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_25/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_30/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_44/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_38/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_13/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_43/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_12/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_22/SL
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_41/SL chip_half_frame_0/gf180mcu_ocd_io__bi_a_35/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_16/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_10/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_40/OE chip_half_frame_0/gf180mcu_ocd_io__bi_a_3/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/A WEN2 chip_half_frame_0/gf180mcu_ocd_io__bi_a_1/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_27/OE ocd_mux_array_1/Y[4] ocd_mux_array_0/Y[6]
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_32/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_11/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_14/IE chip_half_frame_0/gf180mcu_ocd_io__bi_a_0/IE
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_4/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_17/A
+ chip_half_frame_0/gf180mcu_ocd_io__bi_a_19/A chip_half_frame_0/gf180mcu_ocd_io__bi_a_24/OE
+ VSS chip_half_frame
.ends

